// pcie_gen2x8_13_0.v

// Generated using ACDS version 13.0 156 at 2013.06.21.16:21:56

`timescale 1 ps / 1 ps
module pcie_gen2x8_13_1 #(

parameter   PORTS                       = 12,
parameter   BALI                        = 0   )

(
    output [69:0]    fc_reconfig_to_xcvr,
	  input  [45:0]    fc_reconfig_from_xcvr,

		input  wire [31:0] iHIP_CTRL_TEST_IN,          //   hip_ctrl.test_in
		input  wire        iHIP_CTRL_SIMU_MODE_PIPE,   //           .simu_mode_pipe
		input wire iRST_100M_N,
		input wire [PORTS-1:0] iRST_PCIE_N,
		input wire             iRST_CHIP_PCIE_N,
  //////////////////////////////////////////////////////////////////////
  // debug status
  //////////////////////////////////////////////////////////////////////
  output [3:0]        oLANE_ACT,
  output [4:0]        oLTSSM,
  output [1:0]        oCURRENT_SPEED,
  output [31:0]       oPCIE_MISC_STATUS,

		input  wire        iHIP_SERIAL_RX_IN0,         // hip_serial.rx_in0
		input  wire        iHIP_SERIAL_RX_IN1,         //           .rx_in1
		input  wire        iHIP_SERIAL_RX_IN2,         //           .rx_in2
		input  wire        iHIP_SERIAL_RX_IN3,         //           .rx_in3
		input  wire        iHIP_SERIAL_RX_IN4,         //           .rx_in4
		input  wire        iHIP_SERIAL_RX_IN5,         //           .rx_in5
		input  wire        iHIP_SERIAL_RX_IN6,         //           .rx_in6
		input  wire        iHIP_SERIAL_RX_IN7,         //           .rx_in7
		output wire        oHIP_SERIAL_TX_OUT0,        //           .tx_out0
		output wire        oHIP_SERIAL_TX_OUT1,        //           .tx_out1
		output wire        oHIP_SERIAL_TX_OUT2,        //           .tx_out2
		output wire        oHIP_SERIAL_TX_OUT3,        //           .tx_out3
		output wire        oHIP_SERIAL_TX_OUT4,        //           .tx_out4
		output wire        oHIP_SERIAL_TX_OUT5,        //           .tx_out5
		output wire        oHIP_SERIAL_TX_OUT6,        //           .tx_out6
		output wire        oHIP_SERIAL_TX_OUT7,        //           .tx_out7
		input  wire        hip_pipe_sim_pipe_pclk_in, //   hip_pipe.sim_pipe_pclk_in
		output wire [1:0]  hip_pipe_sim_pipe_rate,    //           .sim_pipe_rate
		output wire [4:0]  hip_pipe_sim_ltssmstate,   //           .sim_ltssmstate
		output wire [2:0]  hip_pipe_eidleinfersel0,   //           .eidleinfersel0
		output wire [2:0]  hip_pipe_eidleinfersel1,   //           .eidleinfersel1
		output wire [2:0]  hip_pipe_eidleinfersel2,   //           .eidleinfersel2
		output wire [2:0]  hip_pipe_eidleinfersel3,   //           .eidleinfersel3
		output wire [2:0]  hip_pipe_eidleinfersel4,   //           .eidleinfersel4
		output wire [2:0]  hip_pipe_eidleinfersel5,   //           .eidleinfersel5
		output wire [2:0]  hip_pipe_eidleinfersel6,   //           .eidleinfersel6
		output wire [2:0]  hip_pipe_eidleinfersel7,   //           .eidleinfersel7
		output wire [1:0]  hip_pipe_powerdown0,       //           .powerdown0
		output wire [1:0]  hip_pipe_powerdown1,       //           .powerdown1
		output wire [1:0]  hip_pipe_powerdown2,       //           .powerdown2
		output wire [1:0]  hip_pipe_powerdown3,       //           .powerdown3
		output wire [1:0]  hip_pipe_powerdown4,       //           .powerdown4
		output wire [1:0]  hip_pipe_powerdown5,       //           .powerdown5
		output wire [1:0]  hip_pipe_powerdown6,       //           .powerdown6
		output wire [1:0]  hip_pipe_powerdown7,       //           .powerdown7
		output wire        hip_pipe_rxpolarity0,      //           .rxpolarity0
		output wire        hip_pipe_rxpolarity1,      //           .rxpolarity1
		output wire        hip_pipe_rxpolarity2,      //           .rxpolarity2
		output wire        hip_pipe_rxpolarity3,      //           .rxpolarity3
		output wire        hip_pipe_rxpolarity4,      //           .rxpolarity4
		output wire        hip_pipe_rxpolarity5,      //           .rxpolarity5
		output wire        hip_pipe_rxpolarity6,      //           .rxpolarity6
		output wire        hip_pipe_rxpolarity7,      //           .rxpolarity7
		output wire        hip_pipe_txcompl0,         //           .txcompl0
		output wire        hip_pipe_txcompl1,         //           .txcompl1
		output wire        hip_pipe_txcompl2,         //           .txcompl2
		output wire        hip_pipe_txcompl3,         //           .txcompl3
		output wire        hip_pipe_txcompl4,         //           .txcompl4
		output wire        hip_pipe_txcompl5,         //           .txcompl5
		output wire        hip_pipe_txcompl6,         //           .txcompl6
		output wire        hip_pipe_txcompl7,         //           .txcompl7
		output wire [7:0]  hip_pipe_txdata0,          //           .txdata0
		output wire [7:0]  hip_pipe_txdata1,          //           .txdata1
		output wire [7:0]  hip_pipe_txdata2,          //           .txdata2
		output wire [7:0]  hip_pipe_txdata3,          //           .txdata3
		output wire [7:0]  hip_pipe_txdata4,          //           .txdata4
		output wire [7:0]  hip_pipe_txdata5,          //           .txdata5
		output wire [7:0]  hip_pipe_txdata6,          //           .txdata6
		output wire [7:0]  hip_pipe_txdata7,          //           .txdata7
		output wire        hip_pipe_txdatak0,         //           .txdatak0
		output wire        hip_pipe_txdatak1,         //           .txdatak1
		output wire        hip_pipe_txdatak2,         //           .txdatak2
		output wire        hip_pipe_txdatak3,         //           .txdatak3
		output wire        hip_pipe_txdatak4,         //           .txdatak4
		output wire        hip_pipe_txdatak5,         //           .txdatak5
		output wire        hip_pipe_txdatak6,         //           .txdatak6
		output wire        hip_pipe_txdatak7,         //           .txdatak7
		output wire        hip_pipe_txdetectrx0,      //           .txdetectrx0
		output wire        hip_pipe_txdetectrx1,      //           .txdetectrx1
		output wire        hip_pipe_txdetectrx2,      //           .txdetectrx2
		output wire        hip_pipe_txdetectrx3,      //           .txdetectrx3
		output wire        hip_pipe_txdetectrx4,      //           .txdetectrx4
		output wire        hip_pipe_txdetectrx5,      //           .txdetectrx5
		output wire        hip_pipe_txdetectrx6,      //           .txdetectrx6
		output wire        hip_pipe_txdetectrx7,      //           .txdetectrx7
		output wire        hip_pipe_txelecidle0,      //           .txelecidle0
		output wire        hip_pipe_txelecidle1,      //           .txelecidle1
		output wire        hip_pipe_txelecidle2,      //           .txelecidle2
		output wire        hip_pipe_txelecidle3,      //           .txelecidle3
		output wire        hip_pipe_txelecidle4,      //           .txelecidle4
		output wire        hip_pipe_txelecidle5,      //           .txelecidle5
		output wire        hip_pipe_txelecidle6,      //           .txelecidle6
		output wire        hip_pipe_txelecidle7,      //           .txelecidle7
		output wire        hip_pipe_txdeemph0,        //           .txdeemph0
		output wire        hip_pipe_txdeemph1,        //           .txdeemph1
		output wire        hip_pipe_txdeemph2,        //           .txdeemph2
		output wire        hip_pipe_txdeemph3,        //           .txdeemph3
		output wire        hip_pipe_txdeemph4,        //           .txdeemph4
		output wire        hip_pipe_txdeemph5,        //           .txdeemph5
		output wire        hip_pipe_txdeemph6,        //           .txdeemph6
		output wire        hip_pipe_txdeemph7,        //           .txdeemph7
		output wire [2:0]  hip_pipe_txmargin0,        //           .txmargin0
		output wire [2:0]  hip_pipe_txmargin1,        //           .txmargin1
		output wire [2:0]  hip_pipe_txmargin2,        //           .txmargin2
		output wire [2:0]  hip_pipe_txmargin3,        //           .txmargin3
		output wire [2:0]  hip_pipe_txmargin4,        //           .txmargin4
		output wire [2:0]  hip_pipe_txmargin5,        //           .txmargin5
		output wire [2:0]  hip_pipe_txmargin6,        //           .txmargin6
		output wire [2:0]  hip_pipe_txmargin7,        //           .txmargin7
		output wire        hip_pipe_txswing0,         //           .txswing0
		output wire        hip_pipe_txswing1,         //           .txswing1
		output wire        hip_pipe_txswing2,         //           .txswing2
		output wire        hip_pipe_txswing3,         //           .txswing3
		output wire        hip_pipe_txswing4,         //           .txswing4
		output wire        hip_pipe_txswing5,         //           .txswing5
		output wire        hip_pipe_txswing6,         //           .txswing6
		output wire        hip_pipe_txswing7,         //           .txswing7
		input  wire        hip_pipe_phystatus0,       //           .phystatus0
		input  wire        hip_pipe_phystatus1,       //           .phystatus1
		input  wire        hip_pipe_phystatus2,       //           .phystatus2
		input  wire        hip_pipe_phystatus3,       //           .phystatus3
		input  wire        hip_pipe_phystatus4,       //           .phystatus4
		input  wire        hip_pipe_phystatus5,       //           .phystatus5
		input  wire        hip_pipe_phystatus6,       //           .phystatus6
		input  wire        hip_pipe_phystatus7,       //           .phystatus7
		input  wire [7:0]  hip_pipe_rxdata0,          //           .rxdata0
		input  wire [7:0]  hip_pipe_rxdata1,          //           .rxdata1
		input  wire [7:0]  hip_pipe_rxdata2,          //           .rxdata2
		input  wire [7:0]  hip_pipe_rxdata3,          //           .rxdata3
		input  wire [7:0]  hip_pipe_rxdata4,          //           .rxdata4
		input  wire [7:0]  hip_pipe_rxdata5,          //           .rxdata5
		input  wire [7:0]  hip_pipe_rxdata6,          //           .rxdata6
		input  wire [7:0]  hip_pipe_rxdata7,          //           .rxdata7
		input  wire        hip_pipe_rxdatak0,         //           .rxdatak0
		input  wire        hip_pipe_rxdatak1,         //           .rxdatak1
		input  wire        hip_pipe_rxdatak2,         //           .rxdatak2
		input  wire        hip_pipe_rxdatak3,         //           .rxdatak3
		input  wire        hip_pipe_rxdatak4,         //           .rxdatak4
		input  wire        hip_pipe_rxdatak5,         //           .rxdatak5
		input  wire        hip_pipe_rxdatak6,         //           .rxdatak6
		input  wire        hip_pipe_rxdatak7,         //           .rxdatak7
		input  wire        hip_pipe_rxelecidle0,      //           .rxelecidle0
		input  wire        hip_pipe_rxelecidle1,      //           .rxelecidle1
		input  wire        hip_pipe_rxelecidle2,      //           .rxelecidle2
		input  wire        hip_pipe_rxelecidle3,      //           .rxelecidle3
		input  wire        hip_pipe_rxelecidle4,      //           .rxelecidle4
		input  wire        hip_pipe_rxelecidle5,      //           .rxelecidle5
		input  wire        hip_pipe_rxelecidle6,      //           .rxelecidle6
		input  wire        hip_pipe_rxelecidle7,      //           .rxelecidle7
		input  wire [2:0]  hip_pipe_rxstatus0,        //           .rxstatus0
		input  wire [2:0]  hip_pipe_rxstatus1,        //           .rxstatus1
		input  wire [2:0]  hip_pipe_rxstatus2,        //           .rxstatus2
		input  wire [2:0]  hip_pipe_rxstatus3,        //           .rxstatus3
		input  wire [2:0]  hip_pipe_rxstatus4,        //           .rxstatus4
		input  wire [2:0]  hip_pipe_rxstatus5,        //           .rxstatus5
		input  wire [2:0]  hip_pipe_rxstatus6,        //           .rxstatus6
		input  wire [2:0]  hip_pipe_rxstatus7,        //           .rxstatus7
		input  wire        hip_pipe_rxvalid0,         //           .rxvalid0
		input  wire        hip_pipe_rxvalid1,         //           .rxvalid1
		input  wire        hip_pipe_rxvalid2,         //           .rxvalid2
		input  wire        hip_pipe_rxvalid3,         //           .rxvalid3
		input  wire        hip_pipe_rxvalid4,         //           .rxvalid4
		input  wire        hip_pipe_rxvalid5,         //           .rxvalid5
		input  wire        hip_pipe_rxvalid6,         //           .rxvalid6
		input  wire        hip_pipe_rxvalid7,         //           .rxvalid7
		input  wire        iREF_CLK,                //     refclk.clk
		input  wire        iRST_NPOR_n,            //  pcie_rstn.npor
		input  wire        iPIN_PERST_n,       //           .pin_perst
		input  wire        iRECONFIG_XCVR_CLK,                   //        clk.clk
		input  wire        reset_reset_n,              //      reset.reset_n
  //////////////////////////////////////////////////////////////////////
  // MM DECODE I/F
  //////////////////////////////////////////////////////////////////////
  output [63:0]       oPCIE2MM_WR_DATA,
  output [20:0]       oPCIE2MM_ADDRESS,
  output              oPCIE2MM_WR_EN,
  output              oPCIE2MM_RD_EN,
  input               iMM2PCIE_ACK,
  input  [63:0]       iMM2PCIE_RD_DATA,
  //////////////////////////////////////////////////////////////////////
  // PCIE MM Register I/F
  //////////////////////////////////////////////////////////////////////
  input  [63:0]       iMM_WR_DATA,
  input  [20:0]       iMM_ADDR,
  input               iMM_WR_EN,
  input               iMM_RD_EN,
  output [63:0]       oMM_RD_DATA,
  output              oMM_RD_DATA_V,
  //////////////////////////////////////////////////////////////////////
  // DMA WRITE to DPL BUFFER I/F
  //////////////////////////////////////////////////////////////////////
  input  [PORTS-1:0]  iDPLBUF_REQ,
  output [PORTS-1:0]  oDPLBUF_GNT,

  input  [255:0]      iDPLBUF_DATA,
  input  [PORTS-1:0]  iDPLBUF_DATA_V,
  output              oAPP_RST_n_STATUS,
  //////////////////////////////////////////////////////////////////////
  // Clocks
  //////////////////////////////////////////////////////////////////////
  output              oCLK_PCIE_CORECLKOUT_HIP,
  input               iCLK_PCIE_GLOBAL,
  input               iCLK_100M


	);

	wire          apps_int_msi_app_msi_req;                               // APPS:app_msi_req -> pcie_gen2x8_inst:app_msi_req
	wire          pcie_gen2x8_inst_int_msi_app_msi_ack;                   // pcie_gen2x8_inst:app_msi_ack -> APPS:app_msi_ack
	wire    [0:0] apps_int_msi_app_int_sts;                               // APPS:app_int_sts -> pcie_gen2x8_inst:app_int_sts
	wire          pcie_gen2x8_inst_int_msi_app_int_ack;                   // pcie_gen2x8_inst:app_int_ack -> APPS:app_int_ack
	wire    [2:0] apps_int_msi_app_msi_tc;                                // APPS:app_msi_tc -> pcie_gen2x8_inst:app_msi_tc
	wire    [4:0] apps_int_msi_app_msi_num;                               // APPS:app_msi_num -> pcie_gen2x8_inst:app_msi_num
	wire          apps_config_tl_cpl_pending;                             // APPS:cpl_pending -> pcie_gen2x8_inst:cpl_pending
	wire   [52:0] pcie_gen2x8_inst_config_tl_tl_cfg_sts;                  // pcie_gen2x8_inst:tl_cfg_sts -> APPS:tl_cfg_sts
	wire   [31:0] pcie_gen2x8_inst_config_tl_tl_cfg_ctl;                  // pcie_gen2x8_inst:tl_cfg_ctl -> APPS:tl_cfg_ctl
	wire    [3:0] pcie_gen2x8_inst_config_tl_tl_cfg_add;                  // pcie_gen2x8_inst:tl_cfg_add -> APPS:tl_cfg_add
	wire    [4:0] apps_config_tl_hpg_ctrler;                              // APPS:hpg_ctrler -> pcie_gen2x8_inst:hpg_ctrler
	wire    [6:0] apps_config_tl_cpl_err;                                 // APPS:cpl_err -> pcie_gen2x8_inst:cpl_err
	wire          pcie_gen2x8_inst_power_mngt_pme_to_sr;                  // pcie_gen2x8_inst:pme_to_sr -> APPS:pme_to_sr
	wire          apps_power_mngt_pm_auxpwr;                              // APPS:pm_auxpwr -> pcie_gen2x8_inst:pm_auxpwr
	wire    [9:0] apps_power_mngt_pm_data;                                // APPS:pm_data -> pcie_gen2x8_inst:pm_data
	wire          apps_power_mngt_pme_to_cr;                              // APPS:pme_to_cr -> pcie_gen2x8_inst:pme_to_cr
	wire          apps_power_mngt_pm_event;                               // APPS:pm_event -> pcie_gen2x8_inst:pm_event
	wire          pcie_gen2x8_inst_hip_status_ev128ns;                    // pcie_gen2x8_inst:ev128ns -> APPS:ev128ns
	wire    [3:0] pcie_gen2x8_inst_hip_status_int_status;                 // pcie_gen2x8_inst:int_status -> APPS:int_status
	wire          pcie_gen2x8_inst_hip_status_ev1us;                      // pcie_gen2x8_inst:ev1us -> APPS:ev1us
	wire          pcie_gen2x8_inst_hip_status_derr_cor_ext_rcv;           // pcie_gen2x8_inst:derr_cor_ext_rcv -> APPS:derr_cor_ext_rcv
	wire    [4:0] pcie_gen2x8_inst_hip_status_ltssmstate;                 // pcie_gen2x8_inst:ltssmstate -> APPS:ltssmstate
	wire          pcie_gen2x8_inst_hip_status_rx_par_err;                 // pcie_gen2x8_inst:rx_par_err -> APPS:rx_par_err
	wire          pcie_gen2x8_inst_hip_status_derr_rpl;                   // pcie_gen2x8_inst:derr_rpl -> APPS:derr_rpl
	wire          pcie_gen2x8_inst_hip_status_l2_exit;                    // pcie_gen2x8_inst:l2_exit -> APPS:l2_exit
	wire          pcie_gen2x8_inst_hip_status_cfg_par_err;                // pcie_gen2x8_inst:cfg_par_err -> APPS:cfg_par_err
	wire    [3:0] pcie_gen2x8_inst_hip_status_lane_act;                   // pcie_gen2x8_inst:lane_act -> APPS:lane_act
	wire          pcie_gen2x8_inst_hip_status_dlup_exit;                  // pcie_gen2x8_inst:dlup_exit -> APPS:dlup_exit
	wire    [7:0] pcie_gen2x8_inst_hip_status_ko_cpl_spc_header;          // pcie_gen2x8_inst:ko_cpl_spc_header -> APPS:ko_cpl_spc_header
	wire          pcie_gen2x8_inst_hip_status_hotrst_exit;                // pcie_gen2x8_inst:hotrst_exit -> APPS:hotrst_exit
	wire   [11:0] pcie_gen2x8_inst_hip_status_ko_cpl_spc_data;            // pcie_gen2x8_inst:ko_cpl_spc_data -> APPS:ko_cpl_spc_data
	wire    [1:0] pcie_gen2x8_inst_hip_status_tx_par_err;                 // pcie_gen2x8_inst:tx_par_err -> APPS:tx_par_err
	wire          pcie_gen2x8_inst_hip_status_dlup;                       // pcie_gen2x8_inst:dlup -> APPS:dlup
	wire          pcie_gen2x8_inst_hip_status_derr_cor_ext_rpl;           // pcie_gen2x8_inst:derr_cor_ext_rpl -> APPS:derr_cor_ext_rpl
	wire   [11:0] pcie_gen2x8_inst_tx_cred_tx_cred_datafccp;              // pcie_gen2x8_inst:tx_cred_datafccp -> APPS:tx_cred_datafccp
	wire    [7:0] pcie_gen2x8_inst_tx_cred_tx_cred_hdrfcnp;               // pcie_gen2x8_inst:tx_cred_hdrfcnp -> APPS:tx_cred_hdrfcnp
	wire    [7:0] pcie_gen2x8_inst_tx_cred_tx_cred_hdrfccp;               // pcie_gen2x8_inst:tx_cred_hdrfccp -> APPS:tx_cred_hdrfccp
	wire    [5:0] pcie_gen2x8_inst_tx_cred_tx_cred_fchipcons;             // pcie_gen2x8_inst:tx_cred_fchipcons -> APPS:tx_cred_fchipcons
	wire    [7:0] pcie_gen2x8_inst_tx_cred_tx_cred_hdrfcp;                // pcie_gen2x8_inst:tx_cred_hdrfcp -> APPS:tx_cred_hdrfcp
	wire   [11:0] pcie_gen2x8_inst_tx_cred_tx_cred_datafcp;               // pcie_gen2x8_inst:tx_cred_datafcp -> APPS:tx_cred_datafcp
	wire    [5:0] pcie_gen2x8_inst_tx_cred_tx_cred_fcinfinite;            // pcie_gen2x8_inst:tx_cred_fcinfinite -> APPS:tx_cred_fcinfinite
	wire   [11:0] pcie_gen2x8_inst_tx_cred_tx_cred_datafcnp;              // pcie_gen2x8_inst:tx_cred_datafcnp -> APPS:tx_cred_datafcnp
	wire          apps_rx_bar_be_rx_st_mask;                              // APPS:rx_st_mask -> pcie_gen2x8_inst:rx_st_mask
	wire   [31:0] pcie_gen2x8_inst_rx_bar_be_rx_st_be;                    // pcie_gen2x8_inst:rx_st_be -> APPS:rx_st_be
	wire    [7:0] pcie_gen2x8_inst_rx_bar_be_rx_st_bar;                   // pcie_gen2x8_inst:rx_st_bar -> APPS:rx_st_bar
	wire    [0:0] apps_tx_st_endofpacket;                                 // APPS:tx_st_eop -> pcie_gen2x8_inst:tx_st_eop
	wire    [0:0] apps_tx_st_valid;                                       // APPS:tx_st_valid -> pcie_gen2x8_inst:tx_st_valid
	wire    [0:0] apps_tx_st_startofpacket;                               // APPS:tx_st_sop -> pcie_gen2x8_inst:tx_st_sop
	wire    [0:0] apps_tx_st_error;                                       // APPS:tx_st_err -> pcie_gen2x8_inst:tx_st_err
	wire  [255:0] apps_tx_st_data;                                        // APPS:tx_st_data -> pcie_gen2x8_inst:tx_st_data
	wire    [1:0] apps_tx_st_empty;                                       // APPS:tx_st_empty -> pcie_gen2x8_inst:tx_st_empty
	wire          apps_tx_st_ready;                                       // pcie_gen2x8_inst:tx_st_ready -> APPS:tx_st_ready
	wire   [31:0] pcie_gen2x8_inst_lmi_lmi_dout;                          // pcie_gen2x8_inst:lmi_dout -> APPS:lmi_dout
	wire          apps_lmi_lmi_wren;                                      // APPS:lmi_wren -> pcie_gen2x8_inst:lmi_wren
	wire   [31:0] apps_lmi_lmi_din;                                       // APPS:lmi_din -> pcie_gen2x8_inst:lmi_din
	wire          apps_lmi_lmi_rden;                                      // APPS:lmi_rden -> pcie_gen2x8_inst:lmi_rden
	wire   [11:0] apps_lmi_lmi_addr;                                      // APPS:lmi_addr -> pcie_gen2x8_inst:lmi_addr
	wire          pcie_gen2x8_inst_lmi_lmi_ack;                           // pcie_gen2x8_inst:lmi_ack -> APPS:lmi_ack
	wire    [0:0] pcie_gen2x8_inst_rx_st_endofpacket;                     // pcie_gen2x8_inst:rx_st_eop -> APPS:rx_st_eop
	wire    [0:0] pcie_gen2x8_inst_rx_st_valid;                           // pcie_gen2x8_inst:rx_st_valid -> APPS:rx_st_valid
	wire    [0:0] pcie_gen2x8_inst_rx_st_startofpacket;                   // pcie_gen2x8_inst:rx_st_sop -> APPS:rx_st_sop
	wire    [0:0] pcie_gen2x8_inst_rx_st_error;                           // pcie_gen2x8_inst:rx_st_err -> APPS:rx_st_err
	wire  [255:0] pcie_gen2x8_inst_rx_st_data;                            // pcie_gen2x8_inst:rx_st_data -> APPS:rx_st_data
	wire    [1:0] pcie_gen2x8_inst_rx_st_empty;                           // pcie_gen2x8_inst:rx_st_empty -> APPS:rx_st_empty
	wire          pcie_gen2x8_inst_rx_st_ready;                           // APPS:rx_st_ready -> pcie_gen2x8_inst:rx_st_ready
	wire          pcie_gen2x8_inst_hip_rst_serdes_pll_locked;             // pcie_gen2x8_inst:serdes_pll_locked -> APPS:serdes_pll_locked
	wire          apps_hip_rst_pld_core_ready;                            // APPS:pld_core_ready -> pcie_gen2x8_inst:pld_core_ready
	wire          pcie_gen2x8_inst_hip_rst_pld_clk_inuse;                 // pcie_gen2x8_inst:pld_clk_inuse -> APPS:pld_clk_inuse
	wire          pcie_gen2x8_inst_hip_rst_reset_status;                  // pcie_gen2x8_inst:reset_status -> APPS:reset_status
	wire          pcie_gen2x8_inst_hip_rst_testin_zero;                   // pcie_gen2x8_inst:testin_zero -> APPS:testin_zero
	wire          pcie_gen2x8_inst_coreclkout_hip_clk;                    // pcie_gen2x8_inst:coreclkout_hip -> APPS:coreclkout_hip
	wire          apps_pld_clk_hip_clk;                                   // APPS:pld_clk_hip -> [pcie_gen2x8_inst:pld_clk, pcie_reconfig_driver_0:pld_clk]
	wire  [769:0] alt_xcvr_reconfig_0_reconfig_to_xcvr_reconfig_to_xcvr;  // alt_xcvr_reconfig_0:reconfig_to_xcvr -> pcie_gen2x8_inst:reconfig_to_xcvr
	wire  [505:0] pcie_gen2x8_inst_reconfig_from_xcvr_reconfig_from_xcvr; // pcie_gen2x8_inst:reconfig_from_xcvr -> alt_xcvr_reconfig_0:reconfig_from_xcvr
	wire          pcie_reconfig_driver_0_reconfig_mgmt_waitrequest;       // alt_xcvr_reconfig_0:reconfig_mgmt_waitrequest -> pcie_reconfig_driver_0:reconfig_mgmt_waitrequest
	wire   [31:0] pcie_reconfig_driver_0_reconfig_mgmt_writedata;         // pcie_reconfig_driver_0:reconfig_mgmt_writedata -> alt_xcvr_reconfig_0:reconfig_mgmt_writedata
	wire    [6:0] pcie_reconfig_driver_0_reconfig_mgmt_address;           // pcie_reconfig_driver_0:reconfig_mgmt_address -> alt_xcvr_reconfig_0:reconfig_mgmt_address
	wire          pcie_reconfig_driver_0_reconfig_mgmt_write;             // pcie_reconfig_driver_0:reconfig_mgmt_write -> alt_xcvr_reconfig_0:reconfig_mgmt_write
	wire          pcie_reconfig_driver_0_reconfig_mgmt_read;              // pcie_reconfig_driver_0:reconfig_mgmt_read -> alt_xcvr_reconfig_0:reconfig_mgmt_read
	wire   [31:0] pcie_reconfig_driver_0_reconfig_mgmt_readdata;          // alt_xcvr_reconfig_0:reconfig_mgmt_readdata -> pcie_reconfig_driver_0:reconfig_mgmt_readdata
	wire    [1:0] pcie_gen2x8_inst_hip_currentspeed_currentspeed;         // pcie_gen2x8_inst:currentspeed -> pcie_reconfig_driver_0:currentspeed
	wire          alt_xcvr_reconfig_0_reconfig_busy_reconfig_busy;        // alt_xcvr_reconfig_0:reconfig_busy -> pcie_reconfig_driver_0:reconfig_busy
	wire          apps_hip_status_drv_ev128ns;                            // APPS:ev128ns_drv -> pcie_reconfig_driver_0:ev128ns_drv
	wire    [3:0] apps_hip_status_drv_int_status;                         // APPS:int_status_drv -> pcie_reconfig_driver_0:int_status_drv
	wire          apps_hip_status_drv_ev1us;                              // APPS:ev1us_drv -> pcie_reconfig_driver_0:ev1us_drv
	wire          apps_hip_status_drv_derr_cor_ext_rcv;                   // APPS:derr_cor_ext_rcv_drv -> pcie_reconfig_driver_0:derr_cor_ext_rcv_drv
	wire    [4:0] apps_hip_status_drv_ltssmstate;                         // APPS:ltssmstate_drv -> pcie_reconfig_driver_0:ltssmstate_drv
	wire          apps_hip_status_drv_rx_par_err;                         // APPS:rx_par_err_drv -> pcie_reconfig_driver_0:rx_par_err_drv
	wire          apps_hip_status_drv_derr_rpl;                           // APPS:derr_rpl_drv -> pcie_reconfig_driver_0:derr_rpl_drv
	wire          apps_hip_status_drv_l2_exit;                            // APPS:l2_exit_drv -> pcie_reconfig_driver_0:l2_exit_drv
	wire          apps_hip_status_drv_cfg_par_err;                        // APPS:cfg_par_err_drv -> pcie_reconfig_driver_0:cfg_par_err_drv
	wire    [3:0] apps_hip_status_drv_lane_act;                           // APPS:lane_act_drv -> pcie_reconfig_driver_0:lane_act_drv
	wire          apps_hip_status_drv_dlup_exit;                          // APPS:dlup_exit_drv -> pcie_reconfig_driver_0:dlup_exit_drv
	wire    [7:0] apps_hip_status_drv_ko_cpl_spc_header;                  // APPS:ko_cpl_spc_header_drv -> pcie_reconfig_driver_0:ko_cpl_spc_header_drv
	wire          apps_hip_status_drv_hotrst_exit;                        // APPS:hotrst_exit_drv -> pcie_reconfig_driver_0:hotrst_exit_drv
	wire   [11:0] apps_hip_status_drv_ko_cpl_spc_data;                    // APPS:ko_cpl_spc_data_drv -> pcie_reconfig_driver_0:ko_cpl_spc_data_drv
	wire    [1:0] apps_hip_status_drv_tx_par_err;                         // APPS:tx_par_err_drv -> pcie_reconfig_driver_0:tx_par_err_drv
	wire          apps_hip_status_drv_dlup;                               // APPS:dlup_drv -> pcie_reconfig_driver_0:dlup_drv
	wire          apps_hip_status_drv_derr_cor_ext_rpl;                   // APPS:derr_cor_ext_rpl_drv -> pcie_reconfig_driver_0:derr_cor_ext_rpl_drv
	wire          rst_controller_reset_out_reset;                         // rst_controller:reset_out -> [alt_xcvr_reconfig_0:mgmt_rst_reset, pcie_reconfig_driver_0:reconfig_xcvr_rst]

	altpcie_sv_hip_ast_hwtcl #(
		.lane_mask_hwtcl                          ("x8"),
		.gen123_lane_rate_mode_hwtcl              ("Gen2 (5.0 Gbps)"),
		.port_type_hwtcl                          ("Native endpoint"),
		.pcie_spec_version_hwtcl                  ("2.1"),
		.ast_width_hwtcl                          ("Avalon-ST 256-bit"),
		.pll_refclk_freq_hwtcl                    ("100 MHz"),
		.set_pld_clk_x1_625MHz_hwtcl              (0),
		.use_ast_parity                           (0),
		.multiple_packets_per_cycle_hwtcl         (0),
		.in_cvp_mode_hwtcl                        (0),
		.use_pci_ext_hwtcl                        (0),
		.use_pcie_ext_hwtcl                       (0),
		.use_config_bypass_hwtcl                  (0),
		.hip_reconfig_hwtcl                       (0),
		.enable_tl_only_sim_hwtcl                 (0),
		.bar0_size_mask_hwtcl                     (0),
		.bar0_io_space_hwtcl                      ("Disabled"),
		.bar0_64bit_mem_space_hwtcl               ("Disabled"),
		.bar0_prefetchable_hwtcl                  ("Disabled"),
		.bar1_size_mask_hwtcl                     (0),
		.bar1_io_space_hwtcl                      ("Disabled"),
		.bar1_prefetchable_hwtcl                  ("Disabled"),
		.bar2_size_mask_hwtcl                     (24),
		.bar2_io_space_hwtcl                      ("Disabled"),
		.bar2_64bit_mem_space_hwtcl               ("Disabled"),
		.bar2_prefetchable_hwtcl                  ("Disabled"),
		.bar3_size_mask_hwtcl                     (0),
		.bar3_io_space_hwtcl                      ("Disabled"),
		.bar3_prefetchable_hwtcl                  ("Disabled"),
		.bar4_size_mask_hwtcl                     (0),
		.bar4_io_space_hwtcl                      ("Disabled"),
		.bar4_64bit_mem_space_hwtcl               ("Disabled"),
		.bar4_prefetchable_hwtcl                  ("Disabled"),
		.bar5_size_mask_hwtcl                     (0),
		.bar5_io_space_hwtcl                      ("Disabled"),
		.bar5_prefetchable_hwtcl                  ("Disabled"),
		.expansion_base_address_register_hwtcl    (0),
		.io_window_addr_width_hwtcl               (0),
		.prefetchable_mem_window_addr_width_hwtcl (0),
		.vendor_id_hwtcl                          (7097),
		.device_id_hwtcl                          (4099),
		.revision_id_hwtcl                        (1),
		.class_code_hwtcl                         (16711680),
		.subsystem_vendor_id_hwtcl                (0),
		.subsystem_device_id_hwtcl                (0),
		.max_payload_size_hwtcl                   (2048),
		.extend_tag_field_hwtcl                   ("32"),
		.completion_timeout_hwtcl                 ("ABCD"),
		.enable_completion_timeout_disable_hwtcl  (1),
		.use_aer_hwtcl                            (1),
		.ecrc_check_capable_hwtcl                 (0),
		.ecrc_gen_capable_hwtcl                   (0),
		.use_crc_forwarding_hwtcl                 (0),
		.port_link_number_hwtcl                   (1),
		.dll_active_report_support_hwtcl          (0),
		.surprise_down_error_support_hwtcl        (0),
		.slotclkcfg_hwtcl                         (1),
		.msi_multi_message_capable_hwtcl          ("4"),
		.msi_64bit_addressing_capable_hwtcl       ("true"),
		.msi_masking_capable_hwtcl                ("false"),
		.msi_support_hwtcl                        ("true"),
		.enable_function_msix_support_hwtcl       (0),
		.msix_table_size_hwtcl                    (0),
		.msix_table_offset_hwtcl                  ("0"),
		.msix_table_bir_hwtcl                     (0),
		.msix_pba_offset_hwtcl                    ("0"),
		.msix_pba_bir_hwtcl                       (0),
		.enable_slot_register_hwtcl               (0),
		.slot_power_scale_hwtcl                   (0),
		.slot_power_limit_hwtcl                   (0),
		.slot_number_hwtcl                        (0),
		.endpoint_l0_latency_hwtcl                (0),
		.endpoint_l1_latency_hwtcl                (0),
		.vsec_id_hwtcl                            (40960),
		.vsec_rev_hwtcl                           (0),
		.millisecond_cycle_count_hwtcl            (124250),
		.port_width_be_hwtcl                      (32),
		.port_width_data_hwtcl                    (256),
		.gen3_dcbal_en_hwtcl                      (1),
		.enable_pipe32_sim_hwtcl                  (0),
		.fixed_preset_on                          (0),
		.bypass_cdc_hwtcl                         ("false"),
		.enable_rx_buffer_checking_hwtcl          ("false"),
		.disable_link_x2_support_hwtcl            ("false"),
		.wrong_device_id_hwtcl                    ("disable"),
		.data_pack_rx_hwtcl                       ("disable"),
		.ltssm_1ms_timeout_hwtcl                  ("disable"),
		.ltssm_freqlocked_check_hwtcl             ("disable"),
		.deskew_comma_hwtcl                       ("skp_eieos_deskw"),
		.device_number_hwtcl                      (0),
		.pipex1_debug_sel_hwtcl                   ("disable"),
		.pclk_out_sel_hwtcl                       ("pclk"),
		.no_soft_reset_hwtcl                      ("false"),
		.maximum_current_hwtcl                    (0),
		.d1_support_hwtcl                         ("false"),
		.d2_support_hwtcl                         ("false"),
		.d0_pme_hwtcl                             ("false"),
		.d1_pme_hwtcl                             ("false"),
		.d2_pme_hwtcl                             ("false"),
		.d3_hot_pme_hwtcl                         ("false"),
		.d3_cold_pme_hwtcl                        ("false"),
		.low_priority_vc_hwtcl                    ("single_vc"),
		.disable_snoop_packet_hwtcl               ("false"),
		.enable_l1_aspm_hwtcl                     ("false"),
		.rx_ei_l0s_hwtcl                          (0),
		.enable_l0s_aspm_hwtcl                    ("false"),
		.aspm_config_management_hwtcl             ("true"),
		.l1_exit_latency_sameclock_hwtcl          (0),
		.l1_exit_latency_diffclock_hwtcl          (0),
		.hot_plug_support_hwtcl                   (0),
		.extended_tag_reset_hwtcl                 ("false"),
		.no_command_completed_hwtcl               ("true"),
		.interrupt_pin_hwtcl                      ("inta"),
		.bridge_port_vga_enable_hwtcl             ("false"),
		.bridge_port_ssid_support_hwtcl           ("false"),
		.ssvid_hwtcl                              (0),
		.ssid_hwtcl                               (0),
		.eie_before_nfts_count_hwtcl              (4),
		.gen2_diffclock_nfts_count_hwtcl          (255),
		.gen2_sameclock_nfts_count_hwtcl          (255),
		.l0_exit_latency_sameclock_hwtcl          (6),
		.l0_exit_latency_diffclock_hwtcl          (6),
		.atomic_op_routing_hwtcl                  ("false"),
		.atomic_op_completer_32bit_hwtcl          ("false"),
		.atomic_op_completer_64bit_hwtcl          ("false"),
		.cas_completer_128bit_hwtcl               ("false"),
		.ltr_mechanism_hwtcl                      ("false"),
		.tph_completer_hwtcl                      ("false"),
		.extended_format_field_hwtcl              ("false"),
		.atomic_malformed_hwtcl                   ("true"),
		.flr_capability_hwtcl                     ("false"),
		.enable_adapter_half_rate_mode_hwtcl      ("false"),
		.vc0_clk_enable_hwtcl                     ("true"),
		.register_pipe_signals_hwtcl              ("false"),
		.skp_os_gen3_count_hwtcl                  (0),
		.tx_cdc_almost_empty_hwtcl                (5),
		.rx_l0s_count_idl_hwtcl                   (0),
		.cdc_dummy_insert_limit_hwtcl             (11),
		.ei_delay_powerdown_count_hwtcl           (10),
		.skp_os_schedule_count_hwtcl              (0),
		.fc_init_timer_hwtcl                      (1024),
		.l01_entry_latency_hwtcl                  (31),
		.flow_control_update_count_hwtcl          (30),
		.flow_control_timeout_count_hwtcl         (200),
		.retry_buffer_last_active_address_hwtcl   (2047),
		.reserved_debug_hwtcl                     (0),
		.bypass_clk_switch_hwtcl                  ("true"),
		.l2_async_logic_hwtcl                     ("disable"),
		.indicator_hwtcl                          (0),
		.diffclock_nfts_count_hwtcl               (128),
		.sameclock_nfts_count_hwtcl               (128),
		.rx_cdc_almost_full_hwtcl                 (12),
		.tx_cdc_almost_full_hwtcl                 (11),
		.credit_buffer_allocation_aux_hwtcl       ("absolute"),
		.vc0_rx_flow_ctrl_posted_header_hwtcl     (16),
		.vc0_rx_flow_ctrl_posted_data_hwtcl       (128),
		.vc0_rx_flow_ctrl_nonposted_header_hwtcl  (16),
		.vc0_rx_flow_ctrl_nonposted_data_hwtcl    (0),
		.vc0_rx_flow_ctrl_compl_header_hwtcl      (0),
		.vc0_rx_flow_ctrl_compl_data_hwtcl        (0),
		.cpl_spc_header_hwtcl                     (172),
		.cpl_spc_data_hwtcl                       (692),
		.gen3_rxfreqlock_counter_hwtcl            (0),
		.gen3_skip_ph2_ph3_hwtcl                  (0),
		.g3_bypass_equlz_hwtcl                    (0),
		.cvp_data_compressed_hwtcl                ("false"),
		.cvp_data_encrypted_hwtcl                 ("false"),
		.cvp_mode_reset_hwtcl                     ("false"),
		.cvp_clk_reset_hwtcl                      ("false"),
		.cseb_cpl_status_during_cvp_hwtcl         ("config_retry_status"),
		.core_clk_sel_hwtcl                       ("pld_clk"),
		.cvp_rate_sel_hwtcl                       ("full_rate"),
		.g3_dis_rx_use_prst_hwtcl                 ("true"),
		.g3_dis_rx_use_prst_ep_hwtcl              ("true"),
		.deemphasis_enable_hwtcl                  ("false"),
		.reconfig_to_xcvr_width                   (700),
		.reconfig_from_xcvr_width                 (460),
		.single_rx_detect_hwtcl                   (0),
		.hip_hard_reset_hwtcl                     (0),
		.hwtcl_override_g2_txvod                  (0),
		.rpre_emph_a_val_hwtcl                    (9),
		.rpre_emph_b_val_hwtcl                    (0),
		.rpre_emph_c_val_hwtcl                    (16),
		.rpre_emph_d_val_hwtcl                    (11),
		.rpre_emph_e_val_hwtcl                    (5),
		.rvod_sel_a_val_hwtcl                     (42),
		.rvod_sel_b_val_hwtcl                     (38),
		.rvod_sel_c_val_hwtcl                     (38),
		.rvod_sel_d_val_hwtcl                     (38),
		.rvod_sel_e_val_hwtcl                     (15),
		.hwtcl_override_g3rxcoef                  (0),
		.gen3_coeff_1_hwtcl                       (7),
		.gen3_coeff_1_sel_hwtcl                   ("preset_1"),
		.gen3_coeff_1_preset_hint_hwtcl           (0),
		.gen3_coeff_1_nxtber_more_ptr_hwtcl       (1),
		.gen3_coeff_1_nxtber_more_hwtcl           ("g3_coeff_1_nxtber_more"),
		.gen3_coeff_1_nxtber_less_ptr_hwtcl       (1),
		.gen3_coeff_1_nxtber_less_hwtcl           ("g3_coeff_1_nxtber_less"),
		.gen3_coeff_1_reqber_hwtcl                (0),
		.gen3_coeff_1_ber_meas_hwtcl              (2),
		.gen3_coeff_2_hwtcl                       (0),
		.gen3_coeff_2_sel_hwtcl                   ("preset_2"),
		.gen3_coeff_2_preset_hint_hwtcl           (0),
		.gen3_coeff_2_nxtber_more_ptr_hwtcl       (0),
		.gen3_coeff_2_nxtber_more_hwtcl           ("g3_coeff_2_nxtber_more"),
		.gen3_coeff_2_nxtber_less_ptr_hwtcl       (0),
		.gen3_coeff_2_nxtber_less_hwtcl           ("g3_coeff_2_nxtber_less"),
		.gen3_coeff_2_reqber_hwtcl                (0),
		.gen3_coeff_2_ber_meas_hwtcl              (0),
		.gen3_coeff_3_hwtcl                       (0),
		.gen3_coeff_3_sel_hwtcl                   ("preset_3"),
		.gen3_coeff_3_preset_hint_hwtcl           (0),
		.gen3_coeff_3_nxtber_more_ptr_hwtcl       (0),
		.gen3_coeff_3_nxtber_more_hwtcl           ("g3_coeff_3_nxtber_more"),
		.gen3_coeff_3_nxtber_less_ptr_hwtcl       (0),
		.gen3_coeff_3_nxtber_less_hwtcl           ("g3_coeff_3_nxtber_less"),
		.gen3_coeff_3_reqber_hwtcl                (0),
		.gen3_coeff_3_ber_meas_hwtcl              (0),
		.gen3_coeff_4_hwtcl                       (0),
		.gen3_coeff_4_sel_hwtcl                   ("preset_4"),
		.gen3_coeff_4_preset_hint_hwtcl           (0),
		.gen3_coeff_4_nxtber_more_ptr_hwtcl       (0),
		.gen3_coeff_4_nxtber_more_hwtcl           ("g3_coeff_4_nxtber_more"),
		.gen3_coeff_4_nxtber_less_ptr_hwtcl       (0),
		.gen3_coeff_4_nxtber_less_hwtcl           ("g3_coeff_4_nxtber_less"),
		.gen3_coeff_4_reqber_hwtcl                (0),
		.gen3_coeff_4_ber_meas_hwtcl              (0),
		.gen3_coeff_5_hwtcl                       (0),
		.gen3_coeff_5_sel_hwtcl                   ("preset_5"),
		.gen3_coeff_5_preset_hint_hwtcl           (0),
		.gen3_coeff_5_nxtber_more_ptr_hwtcl       (0),
		.gen3_coeff_5_nxtber_more_hwtcl           ("g3_coeff_5_nxtber_more"),
		.gen3_coeff_5_nxtber_less_ptr_hwtcl       (0),
		.gen3_coeff_5_nxtber_less_hwtcl           ("g3_coeff_5_nxtber_less"),
		.gen3_coeff_5_reqber_hwtcl                (0),
		.gen3_coeff_5_ber_meas_hwtcl              (0),
		.gen3_coeff_6_hwtcl                       (0),
		.gen3_coeff_6_sel_hwtcl                   ("preset_6"),
		.gen3_coeff_6_preset_hint_hwtcl           (0),
		.gen3_coeff_6_nxtber_more_ptr_hwtcl       (0),
		.gen3_coeff_6_nxtber_more_hwtcl           ("g3_coeff_6_nxtber_more"),
		.gen3_coeff_6_nxtber_less_ptr_hwtcl       (0),
		.gen3_coeff_6_nxtber_less_hwtcl           ("g3_coeff_6_nxtber_less"),
		.gen3_coeff_6_reqber_hwtcl                (0),
		.gen3_coeff_6_ber_meas_hwtcl              (0),
		.gen3_coeff_7_hwtcl                       (0),
		.gen3_coeff_7_sel_hwtcl                   ("preset_7"),
		.gen3_coeff_7_preset_hint_hwtcl           (0),
		.gen3_coeff_7_nxtber_more_ptr_hwtcl       (0),
		.gen3_coeff_7_nxtber_more_hwtcl           ("g3_coeff_7_nxtber_more"),
		.gen3_coeff_7_nxtber_less_ptr_hwtcl       (0),
		.gen3_coeff_7_nxtber_less_hwtcl           ("g3_coeff_7_nxtber_less"),
		.gen3_coeff_7_reqber_hwtcl                (0),
		.gen3_coeff_7_ber_meas_hwtcl              (0),
		.gen3_coeff_8_hwtcl                       (0),
		.gen3_coeff_8_sel_hwtcl                   ("preset_8"),
		.gen3_coeff_8_preset_hint_hwtcl           (0),
		.gen3_coeff_8_nxtber_more_ptr_hwtcl       (0),
		.gen3_coeff_8_nxtber_more_hwtcl           ("g3_coeff_8_nxtber_more"),
		.gen3_coeff_8_nxtber_less_ptr_hwtcl       (0),
		.gen3_coeff_8_nxtber_less_hwtcl           ("g3_coeff_8_nxtber_less"),
		.gen3_coeff_8_reqber_hwtcl                (0),
		.gen3_coeff_8_ber_meas_hwtcl              (0),
		.gen3_coeff_9_hwtcl                       (0),
		.gen3_coeff_9_sel_hwtcl                   ("preset_9"),
		.gen3_coeff_9_preset_hint_hwtcl           (0),
		.gen3_coeff_9_nxtber_more_ptr_hwtcl       (0),
		.gen3_coeff_9_nxtber_more_hwtcl           ("g3_coeff_9_nxtber_more"),
		.gen3_coeff_9_nxtber_less_ptr_hwtcl       (0),
		.gen3_coeff_9_nxtber_less_hwtcl           ("g3_coeff_9_nxtber_less"),
		.gen3_coeff_9_reqber_hwtcl                (0),
		.gen3_coeff_9_ber_meas_hwtcl              (0),
		.gen3_coeff_10_hwtcl                      (0),
		.gen3_coeff_10_sel_hwtcl                  ("preset_10"),
		.gen3_coeff_10_preset_hint_hwtcl          (0),
		.gen3_coeff_10_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_10_nxtber_more_hwtcl          ("g3_coeff_10_nxtber_more"),
		.gen3_coeff_10_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_10_nxtber_less_hwtcl          ("g3_coeff_10_nxtber_less"),
		.gen3_coeff_10_reqber_hwtcl               (0),
		.gen3_coeff_10_ber_meas_hwtcl             (0),
		.gen3_coeff_11_hwtcl                      (0),
		.gen3_coeff_11_sel_hwtcl                  ("preset_11"),
		.gen3_coeff_11_preset_hint_hwtcl          (0),
		.gen3_coeff_11_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_11_nxtber_more_hwtcl          ("g3_coeff_11_nxtber_more"),
		.gen3_coeff_11_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_11_nxtber_less_hwtcl          ("g3_coeff_11_nxtber_less"),
		.gen3_coeff_11_reqber_hwtcl               (0),
		.gen3_coeff_11_ber_meas_hwtcl             (0),
		.gen3_coeff_12_hwtcl                      (0),
		.gen3_coeff_12_sel_hwtcl                  ("preset_12"),
		.gen3_coeff_12_preset_hint_hwtcl          (0),
		.gen3_coeff_12_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_12_nxtber_more_hwtcl          ("g3_coeff_12_nxtber_more"),
		.gen3_coeff_12_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_12_nxtber_less_hwtcl          ("g3_coeff_12_nxtber_less"),
		.gen3_coeff_12_reqber_hwtcl               (0),
		.gen3_coeff_12_ber_meas_hwtcl             (0),
		.gen3_coeff_13_hwtcl                      (0),
		.gen3_coeff_13_sel_hwtcl                  ("preset_13"),
		.gen3_coeff_13_preset_hint_hwtcl          (0),
		.gen3_coeff_13_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_13_nxtber_more_hwtcl          ("g3_coeff_13_nxtber_more"),
		.gen3_coeff_13_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_13_nxtber_less_hwtcl          ("g3_coeff_13_nxtber_less"),
		.gen3_coeff_13_reqber_hwtcl               (0),
		.gen3_coeff_13_ber_meas_hwtcl             (0),
		.gen3_coeff_14_hwtcl                      (0),
		.gen3_coeff_14_sel_hwtcl                  ("preset_14"),
		.gen3_coeff_14_preset_hint_hwtcl          (0),
		.gen3_coeff_14_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_14_nxtber_more_hwtcl          ("g3_coeff_14_nxtber_more"),
		.gen3_coeff_14_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_14_nxtber_less_hwtcl          ("g3_coeff_14_nxtber_less"),
		.gen3_coeff_14_reqber_hwtcl               (0),
		.gen3_coeff_14_ber_meas_hwtcl             (0),
		.gen3_coeff_15_hwtcl                      (0),
		.gen3_coeff_15_sel_hwtcl                  ("preset_15"),
		.gen3_coeff_15_preset_hint_hwtcl          (0),
		.gen3_coeff_15_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_15_nxtber_more_hwtcl          ("g3_coeff_15_nxtber_more"),
		.gen3_coeff_15_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_15_nxtber_less_hwtcl          ("g3_coeff_15_nxtber_less"),
		.gen3_coeff_15_reqber_hwtcl               (0),
		.gen3_coeff_15_ber_meas_hwtcl             (0),
		.gen3_coeff_16_hwtcl                      (0),
		.gen3_coeff_16_sel_hwtcl                  ("preset_16"),
		.gen3_coeff_16_preset_hint_hwtcl          (0),
		.gen3_coeff_16_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_16_nxtber_more_hwtcl          ("g3_coeff_16_nxtber_more"),
		.gen3_coeff_16_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_16_nxtber_less_hwtcl          ("g3_coeff_16_nxtber_less"),
		.gen3_coeff_16_reqber_hwtcl               (0),
		.gen3_coeff_16_ber_meas_hwtcl             (0),
		.gen3_coeff_17_hwtcl                      (0),
		.gen3_coeff_17_sel_hwtcl                  ("preset_17"),
		.gen3_coeff_17_preset_hint_hwtcl          (0),
		.gen3_coeff_17_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_17_nxtber_more_hwtcl          ("g3_coeff_17_nxtber_more"),
		.gen3_coeff_17_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_17_nxtber_less_hwtcl          ("g3_coeff_17_nxtber_less"),
		.gen3_coeff_17_reqber_hwtcl               (0),
		.gen3_coeff_17_ber_meas_hwtcl             (0),
		.gen3_coeff_18_hwtcl                      (0),
		.gen3_coeff_18_sel_hwtcl                  ("preset_18"),
		.gen3_coeff_18_preset_hint_hwtcl          (0),
		.gen3_coeff_18_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_18_nxtber_more_hwtcl          ("g3_coeff_18_nxtber_more"),
		.gen3_coeff_18_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_18_nxtber_less_hwtcl          ("g3_coeff_18_nxtber_less"),
		.gen3_coeff_18_reqber_hwtcl               (0),
		.gen3_coeff_18_ber_meas_hwtcl             (0),
		.gen3_coeff_19_hwtcl                      (0),
		.gen3_coeff_19_sel_hwtcl                  ("preset_19"),
		.gen3_coeff_19_preset_hint_hwtcl          (0),
		.gen3_coeff_19_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_19_nxtber_more_hwtcl          ("g3_coeff_19_nxtber_more"),
		.gen3_coeff_19_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_19_nxtber_less_hwtcl          ("g3_coeff_19_nxtber_less"),
		.gen3_coeff_19_reqber_hwtcl               (0),
		.gen3_coeff_19_ber_meas_hwtcl             (0),
		.gen3_coeff_20_hwtcl                      (0),
		.gen3_coeff_20_sel_hwtcl                  ("preset_20"),
		.gen3_coeff_20_preset_hint_hwtcl          (0),
		.gen3_coeff_20_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_20_nxtber_more_hwtcl          ("g3_coeff_20_nxtber_more"),
		.gen3_coeff_20_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_20_nxtber_less_hwtcl          ("g3_coeff_20_nxtber_less"),
		.gen3_coeff_20_reqber_hwtcl               (0),
		.gen3_coeff_20_ber_meas_hwtcl             (0),
		.gen3_coeff_21_hwtcl                      (0),
		.gen3_coeff_21_sel_hwtcl                  ("preset_21"),
		.gen3_coeff_21_preset_hint_hwtcl          (0),
		.gen3_coeff_21_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_21_nxtber_more_hwtcl          ("g3_coeff_21_nxtber_more"),
		.gen3_coeff_21_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_21_nxtber_less_hwtcl          ("g3_coeff_21_nxtber_less"),
		.gen3_coeff_21_reqber_hwtcl               (0),
		.gen3_coeff_21_ber_meas_hwtcl             (0),
		.gen3_coeff_22_hwtcl                      (0),
		.gen3_coeff_22_sel_hwtcl                  ("preset_22"),
		.gen3_coeff_22_preset_hint_hwtcl          (0),
		.gen3_coeff_22_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_22_nxtber_more_hwtcl          ("g3_coeff_22_nxtber_more"),
		.gen3_coeff_22_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_22_nxtber_less_hwtcl          ("g3_coeff_22_nxtber_less"),
		.gen3_coeff_22_reqber_hwtcl               (0),
		.gen3_coeff_22_ber_meas_hwtcl             (0),
		.gen3_coeff_23_hwtcl                      (0),
		.gen3_coeff_23_sel_hwtcl                  ("preset_23"),
		.gen3_coeff_23_preset_hint_hwtcl          (0),
		.gen3_coeff_23_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_23_nxtber_more_hwtcl          ("g3_coeff_23_nxtber_more"),
		.gen3_coeff_23_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_23_nxtber_less_hwtcl          ("g3_coeff_23_nxtber_less"),
		.gen3_coeff_23_reqber_hwtcl               (0),
		.gen3_coeff_23_ber_meas_hwtcl             (0),
		.gen3_coeff_24_hwtcl                      (0),
		.gen3_coeff_24_sel_hwtcl                  ("preset_24"),
		.gen3_coeff_24_preset_hint_hwtcl          (0),
		.gen3_coeff_24_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_24_nxtber_more_hwtcl          ("g3_coeff_24_nxtber_more"),
		.gen3_coeff_24_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_24_nxtber_less_hwtcl          ("g3_coeff_24_nxtber_less"),
		.gen3_coeff_24_reqber_hwtcl               (0),
		.gen3_coeff_24_ber_meas_hwtcl             (0),
		.hwtcl_override_g3txcoef                  (0),
		.gen3_preset_coeff_1_hwtcl                (0),
		.gen3_preset_coeff_2_hwtcl                (0),
		.gen3_preset_coeff_3_hwtcl                (0),
		.gen3_preset_coeff_4_hwtcl                (0),
		.gen3_preset_coeff_5_hwtcl                (0),
		.gen3_preset_coeff_6_hwtcl                (0),
		.gen3_preset_coeff_7_hwtcl                (0),
		.gen3_preset_coeff_8_hwtcl                (0),
		.gen3_preset_coeff_9_hwtcl                (0),
		.gen3_preset_coeff_10_hwtcl               (0),
		.gen3_preset_coeff_11_hwtcl               (0),
		.gen3_low_freq_hwtcl                      (0),
		.full_swing_hwtcl                         (53),
		.gen3_full_swing_hwtcl                    (35),
		.use_atx_pll_hwtcl                        (0),
		.low_latency_mode_hwtcl                   (0)
	) pcie_gen2x8_inst (
		//lz try different reset  .npor                   (iRST_NPOR_n),    //               npor.npor
		.npor                   (iPIN_PERST_n),    //               npor.npor
		.pin_perst              (iPIN_PERST_n),       //                   .pin_perst
		.lmi_addr               (apps_lmi_lmi_addr), //                lmi.lmi_addr
		.lmi_din                (apps_lmi_lmi_din),  //                   .lmi_din
		.lmi_rden               (apps_lmi_lmi_rden), //                   .lmi_rden
		.lmi_wren               (apps_lmi_lmi_wren), //                   .lmi_wren
		.lmi_ack                (pcie_gen2x8_inst_lmi_lmi_ack),          //                   .lmi_ack
		.lmi_dout               (pcie_gen2x8_inst_lmi_lmi_dout),         //                   .lmi_dout
		.hpg_ctrler             (apps_config_tl_hpg_ctrler), //          config_tl.hpg_ctrler
		.tl_cfg_add             (pcie_gen2x8_inst_config_tl_tl_cfg_add), //                   .tl_cfg_add
		.tl_cfg_ctl             (pcie_gen2x8_inst_config_tl_tl_cfg_ctl), //                   .tl_cfg_ctl
		.tl_cfg_sts             (pcie_gen2x8_inst_config_tl_tl_cfg_sts), //                   .tl_cfg_sts
		.cpl_err                (apps_config_tl_cpl_err),    //                   .cpl_err
		.cpl_pending            (apps_config_tl_cpl_pending),//                   .cpl_pending
		.pm_auxpwr              (apps_power_mngt_pm_auxpwr), //         power_mngt.pm_auxpwr
		.pm_data                (apps_power_mngt_pm_data),   //                   .pm_data
		.pme_to_cr              (apps_power_mngt_pme_to_cr), //                   .pme_to_cr
		.pm_event               (apps_power_mngt_pm_event),  //                   .pm_event
		.pme_to_sr              (pcie_gen2x8_inst_power_mngt_pme_to_sr), //                   .pme_to_sr
		.rx_st_sop              (pcie_gen2x8_inst_rx_st_startofpacket),  //              rx_st.startofpacket
		.rx_st_eop              (pcie_gen2x8_inst_rx_st_endofpacket),    //                   .endofpacket
		.rx_st_err              (pcie_gen2x8_inst_rx_st_error),          //                   .error
		.rx_st_valid            (pcie_gen2x8_inst_rx_st_valid),          //                   .valid
		.rx_st_empty            (pcie_gen2x8_inst_rx_st_empty),          //                   .empty
		.rx_st_ready            (pcie_gen2x8_inst_rx_st_ready),          //                   .ready
		.rx_st_data             (pcie_gen2x8_inst_rx_st_data),           //                   .data
		.rx_st_bar              (pcie_gen2x8_inst_rx_bar_be_rx_st_bar),  //          rx_bar_be.rx_st_bar
		.rx_st_be               (pcie_gen2x8_inst_rx_bar_be_rx_st_be),   //                   .rx_st_be
		.rx_st_mask             (apps_rx_bar_be_rx_st_mask), //                   .rx_st_mask
		.tx_st_sop              (apps_tx_st_startofpacket),  //              tx_st.startofpacket
		.tx_st_eop              (apps_tx_st_endofpacket),    //                   .endofpacket
		.tx_st_err              (apps_tx_st_error),  //                   .error
		.tx_st_valid            (apps_tx_st_valid),  //                   .valid
		.tx_st_empty            (apps_tx_st_empty),  //                   .empty
		.tx_st_ready            (apps_tx_st_ready),  //                   .ready
		.tx_st_data             (apps_tx_st_data),   //                   .data
		.tx_cred_datafccp       (pcie_gen2x8_inst_tx_cred_tx_cred_datafccp),     //            tx_cred.tx_cred_datafccp
		.tx_cred_datafcnp       (pcie_gen2x8_inst_tx_cred_tx_cred_datafcnp),     //                   .tx_cred_datafcnp
		.tx_cred_datafcp        (pcie_gen2x8_inst_tx_cred_tx_cred_datafcp),      //                   .tx_cred_datafcp
		.tx_cred_fchipcons      (pcie_gen2x8_inst_tx_cred_tx_cred_fchipcons),    //                   .tx_cred_fchipcons
		.tx_cred_fcinfinite     (pcie_gen2x8_inst_tx_cred_tx_cred_fcinfinite),   //                   .tx_cred_fcinfinite
		.tx_cred_hdrfccp        (pcie_gen2x8_inst_tx_cred_tx_cred_hdrfccp),      //                   .tx_cred_hdrfccp
		.tx_cred_hdrfcnp        (pcie_gen2x8_inst_tx_cred_tx_cred_hdrfcnp),      //                   .tx_cred_hdrfcnp
		.tx_cred_hdrfcp         (pcie_gen2x8_inst_tx_cred_tx_cred_hdrfcp),       //                   .tx_cred_hdrfcp
		.pld_clk                (iCLK_PCIE_GLOBAL),      //            pld_clk.clk
		.coreclkout_hip         (oCLK_PCIE_CORECLKOUT_HIP),   //     coreclkout_hip.clk
		.refclk                 (iREF_CLK),        //             refclk.clk
		.reset_status           (pcie_gen2x8_inst_hip_rst_reset_status), //            hip_rst.reset_status
		.serdes_pll_locked      (pcie_gen2x8_inst_hip_rst_serdes_pll_locked),    //                   .serdes_pll_locked
		.pld_clk_inuse          (pcie_gen2x8_inst_hip_rst_pld_clk_inuse),//                   .pld_clk_inuse
		.pld_core_ready         (apps_hip_rst_pld_core_ready),           //                   .pld_core_ready
		.testin_zero            (pcie_gen2x8_inst_hip_rst_testin_zero),  //                   .testin_zero
		.reconfig_to_xcvr       (alt_xcvr_reconfig_0_reconfig_to_xcvr_reconfig_to_xcvr),  //   reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr     (pcie_gen2x8_inst_reconfig_from_xcvr_reconfig_from_xcvr), // reconfig_from_xcvr.reconfig_from_xcvr
		.rx_in0                 (iHIP_SERIAL_RX_IN0), //         hip_serial.rx_in0
		.rx_in1                 (iHIP_SERIAL_RX_IN1), //                   .rx_in1
		.rx_in2                 (iHIP_SERIAL_RX_IN2), //                   .rx_in2
		.rx_in3                 (iHIP_SERIAL_RX_IN3), //                   .rx_in3
		.rx_in4                 (iHIP_SERIAL_RX_IN4), //                   .rx_in4
		.rx_in5                 (iHIP_SERIAL_RX_IN5), //                   .rx_in5
		.rx_in6                 (iHIP_SERIAL_RX_IN6), //                   .rx_in6
		.rx_in7                 (iHIP_SERIAL_RX_IN7), //                   .rx_in7
		.tx_out0                (oHIP_SERIAL_TX_OUT0),//                   .tx_out0
		.tx_out1                (oHIP_SERIAL_TX_OUT1),//                   .tx_out1
		.tx_out2                (oHIP_SERIAL_TX_OUT2),//                   .tx_out2
		.tx_out3                (oHIP_SERIAL_TX_OUT3),//                   .tx_out3
		.tx_out4                (oHIP_SERIAL_TX_OUT4),//                   .tx_out4
		.tx_out5                (oHIP_SERIAL_TX_OUT5),//                   .tx_out5
		.tx_out6                (oHIP_SERIAL_TX_OUT6),//                   .tx_out6
		.tx_out7                (oHIP_SERIAL_TX_OUT7),//                   .tx_out7
		.sim_pipe_pclk_in       (hip_pipe_sim_pipe_pclk_in), //           hip_pipe.sim_pipe_pclk_in
		.sim_pipe_rate          (hip_pipe_sim_pipe_rate),    //                   .sim_pipe_rate
		.sim_ltssmstate         (hip_pipe_sim_ltssmstate),   //                   .sim_ltssmstate
		.eidleinfersel0         (hip_pipe_eidleinfersel0),   //                   .eidleinfersel0
		.eidleinfersel1         (hip_pipe_eidleinfersel1),   //                   .eidleinfersel1
		.eidleinfersel2         (hip_pipe_eidleinfersel2),   //                   .eidleinfersel2
		.eidleinfersel3         (hip_pipe_eidleinfersel3),   //                   .eidleinfersel3
		.eidleinfersel4         (hip_pipe_eidleinfersel4),   //                   .eidleinfersel4
		.eidleinfersel5         (hip_pipe_eidleinfersel5),   //                   .eidleinfersel5
		.eidleinfersel6         (hip_pipe_eidleinfersel6),   //                   .eidleinfersel6
		.eidleinfersel7         (hip_pipe_eidleinfersel7),   //                   .eidleinfersel7
		.powerdown0             (hip_pipe_powerdown0),       //                   .powerdown0
		.powerdown1             (hip_pipe_powerdown1),       //                   .powerdown1
		.powerdown2             (hip_pipe_powerdown2),       //                   .powerdown2
		.powerdown3             (hip_pipe_powerdown3),       //                   .powerdown3
		.powerdown4             (hip_pipe_powerdown4),       //                   .powerdown4
		.powerdown5             (hip_pipe_powerdown5),       //                   .powerdown5
		.powerdown6             (hip_pipe_powerdown6),       //                   .powerdown6
		.powerdown7             (hip_pipe_powerdown7),       //                   .powerdown7
		.rxpolarity0            (hip_pipe_rxpolarity0),      //                   .rxpolarity0
		.rxpolarity1            (hip_pipe_rxpolarity1),      //                   .rxpolarity1
		.rxpolarity2            (hip_pipe_rxpolarity2),      //                   .rxpolarity2
		.rxpolarity3            (hip_pipe_rxpolarity3),      //                   .rxpolarity3
		.rxpolarity4            (hip_pipe_rxpolarity4),      //                   .rxpolarity4
		.rxpolarity5            (hip_pipe_rxpolarity5),      //                   .rxpolarity5
		.rxpolarity6            (hip_pipe_rxpolarity6),      //                   .rxpolarity6
		.rxpolarity7            (hip_pipe_rxpolarity7),      //                   .rxpolarity7
		.txcompl0               (hip_pipe_txcompl0), //                   .txcompl0
		.txcompl1               (hip_pipe_txcompl1), //                   .txcompl1
		.txcompl2               (hip_pipe_txcompl2), //                   .txcompl2
		.txcompl3               (hip_pipe_txcompl3), //                   .txcompl3
		.txcompl4               (hip_pipe_txcompl4), //                   .txcompl4
		.txcompl5               (hip_pipe_txcompl5), //                   .txcompl5
		.txcompl6               (hip_pipe_txcompl6), //                   .txcompl6
		.txcompl7               (hip_pipe_txcompl7), //                   .txcompl7
		.txdata0                (hip_pipe_txdata0),  //                   .txdata0
		.txdata1                (hip_pipe_txdata1),  //                   .txdata1
		.txdata2                (hip_pipe_txdata2),  //                   .txdata2
		.txdata3                (hip_pipe_txdata3),  //                   .txdata3
		.txdata4                (hip_pipe_txdata4),  //                   .txdata4
		.txdata5                (hip_pipe_txdata5),  //                   .txdata5
		.txdata6                (hip_pipe_txdata6),  //                   .txdata6
		.txdata7                (hip_pipe_txdata7),  //                   .txdata7
		.txdatak0               (hip_pipe_txdatak0), //                   .txdatak0
		.txdatak1               (hip_pipe_txdatak1), //                   .txdatak1
		.txdatak2               (hip_pipe_txdatak2), //                   .txdatak2
		.txdatak3               (hip_pipe_txdatak3), //                   .txdatak3
		.txdatak4               (hip_pipe_txdatak4), //                   .txdatak4
		.txdatak5               (hip_pipe_txdatak5), //                   .txdatak5
		.txdatak6               (hip_pipe_txdatak6), //                   .txdatak6
		.txdatak7               (hip_pipe_txdatak7), //                   .txdatak7
		.txdetectrx0            (hip_pipe_txdetectrx0),      //                   .txdetectrx0
		.txdetectrx1            (hip_pipe_txdetectrx1),      //                   .txdetectrx1
		.txdetectrx2            (hip_pipe_txdetectrx2),      //                   .txdetectrx2
		.txdetectrx3            (hip_pipe_txdetectrx3),      //                   .txdetectrx3
		.txdetectrx4            (hip_pipe_txdetectrx4),      //                   .txdetectrx4
		.txdetectrx5            (hip_pipe_txdetectrx5),      //                   .txdetectrx5
		.txdetectrx6            (hip_pipe_txdetectrx6),      //                   .txdetectrx6
		.txdetectrx7            (hip_pipe_txdetectrx7),      //                   .txdetectrx7
		.txelecidle0            (hip_pipe_txelecidle0),      //                   .txelecidle0
		.txelecidle1            (hip_pipe_txelecidle1),      //                   .txelecidle1
		.txelecidle2            (hip_pipe_txelecidle2),      //                   .txelecidle2
		.txelecidle3            (hip_pipe_txelecidle3),      //                   .txelecidle3
		.txelecidle4            (hip_pipe_txelecidle4),      //                   .txelecidle4
		.txelecidle5            (hip_pipe_txelecidle5),      //                   .txelecidle5
		.txelecidle6            (hip_pipe_txelecidle6),      //                   .txelecidle6
		.txelecidle7            (hip_pipe_txelecidle7),      //                   .txelecidle7
		.txdeemph0              (hip_pipe_txdeemph0),//                   .txdeemph0
		.txdeemph1              (hip_pipe_txdeemph1),//                   .txdeemph1
		.txdeemph2              (hip_pipe_txdeemph2),//                   .txdeemph2
		.txdeemph3              (hip_pipe_txdeemph3),//                   .txdeemph3
		.txdeemph4              (hip_pipe_txdeemph4),//                   .txdeemph4
		.txdeemph5              (hip_pipe_txdeemph5),//                   .txdeemph5
		.txdeemph6              (hip_pipe_txdeemph6),//                   .txdeemph6
		.txdeemph7              (hip_pipe_txdeemph7),//                   .txdeemph7
		.txmargin0              (hip_pipe_txmargin0),//                   .txmargin0
		.txmargin1              (hip_pipe_txmargin1),//                   .txmargin1
		.txmargin2              (hip_pipe_txmargin2),//                   .txmargin2
		.txmargin3              (hip_pipe_txmargin3),//                   .txmargin3
		.txmargin4              (hip_pipe_txmargin4),//                   .txmargin4
		.txmargin5              (hip_pipe_txmargin5),//                   .txmargin5
		.txmargin6              (hip_pipe_txmargin6),//                   .txmargin6
		.txmargin7              (hip_pipe_txmargin7),//                   .txmargin7
		.txswing0               (hip_pipe_txswing0), //                   .txswing0
		.txswing1               (hip_pipe_txswing1), //                   .txswing1
		.txswing2               (hip_pipe_txswing2), //                   .txswing2
		.txswing3               (hip_pipe_txswing3), //                   .txswing3
		.txswing4               (hip_pipe_txswing4), //                   .txswing4
		.txswing5               (hip_pipe_txswing5), //                   .txswing5
		.txswing6               (hip_pipe_txswing6), //                   .txswing6
		.txswing7               (hip_pipe_txswing7), //                   .txswing7
		.phystatus0             (hip_pipe_phystatus0),       //                   .phystatus0
		.phystatus1             (hip_pipe_phystatus1),       //                   .phystatus1
		.phystatus2             (hip_pipe_phystatus2),       //                   .phystatus2
		.phystatus3             (hip_pipe_phystatus3),       //                   .phystatus3
		.phystatus4             (hip_pipe_phystatus4),       //                   .phystatus4
		.phystatus5             (hip_pipe_phystatus5),       //                   .phystatus5
		.phystatus6             (hip_pipe_phystatus6),       //                   .phystatus6
		.phystatus7             (hip_pipe_phystatus7),       //                   .phystatus7
		.rxdata0                (hip_pipe_rxdata0),  //                   .rxdata0
		.rxdata1                (hip_pipe_rxdata1),  //                   .rxdata1
		.rxdata2                (hip_pipe_rxdata2),  //                   .rxdata2
		.rxdata3                (hip_pipe_rxdata3),  //                   .rxdata3
		.rxdata4                (hip_pipe_rxdata4),  //                   .rxdata4
		.rxdata5                (hip_pipe_rxdata5),  //                   .rxdata5
		.rxdata6                (hip_pipe_rxdata6),  //                   .rxdata6
		.rxdata7                (hip_pipe_rxdata7),  //                   .rxdata7
		.rxdatak0               (hip_pipe_rxdatak0), //                   .rxdatak0
		.rxdatak1               (hip_pipe_rxdatak1), //                   .rxdatak1
		.rxdatak2               (hip_pipe_rxdatak2), //                   .rxdatak2
		.rxdatak3               (hip_pipe_rxdatak3), //                   .rxdatak3
		.rxdatak4               (hip_pipe_rxdatak4), //                   .rxdatak4
		.rxdatak5               (hip_pipe_rxdatak5), //                   .rxdatak5
		.rxdatak6               (hip_pipe_rxdatak6), //                   .rxdatak6
		.rxdatak7               (hip_pipe_rxdatak7), //                   .rxdatak7
		.rxelecidle0            (hip_pipe_rxelecidle0),      //                   .rxelecidle0
		.rxelecidle1            (hip_pipe_rxelecidle1),      //                   .rxelecidle1
		.rxelecidle2            (hip_pipe_rxelecidle2),      //                   .rxelecidle2
		.rxelecidle3            (hip_pipe_rxelecidle3),      //                   .rxelecidle3
		.rxelecidle4            (hip_pipe_rxelecidle4),      //                   .rxelecidle4
		.rxelecidle5            (hip_pipe_rxelecidle5),      //                   .rxelecidle5
		.rxelecidle6            (hip_pipe_rxelecidle6),      //                   .rxelecidle6
		.rxelecidle7            (hip_pipe_rxelecidle7),      //                   .rxelecidle7
		.rxstatus0              (hip_pipe_rxstatus0),//                   .rxstatus0
		.rxstatus1              (hip_pipe_rxstatus1),//                   .rxstatus1
		.rxstatus2              (hip_pipe_rxstatus2),//                   .rxstatus2
		.rxstatus3              (hip_pipe_rxstatus3),//                   .rxstatus3
		.rxstatus4              (hip_pipe_rxstatus4),//                   .rxstatus4
		.rxstatus5              (hip_pipe_rxstatus5),//                   .rxstatus5
		.rxstatus6              (hip_pipe_rxstatus6),//                   .rxstatus6
		.rxstatus7              (hip_pipe_rxstatus7),//                   .rxstatus7
		.rxvalid0               (hip_pipe_rxvalid0), //                   .rxvalid0
		.rxvalid1               (hip_pipe_rxvalid1), //                   .rxvalid1
		.rxvalid2               (hip_pipe_rxvalid2), //                   .rxvalid2
		.rxvalid3               (hip_pipe_rxvalid3), //                   .rxvalid3
		.rxvalid4               (hip_pipe_rxvalid4), //                   .rxvalid4
		.rxvalid5               (hip_pipe_rxvalid5), //                   .rxvalid5
		.rxvalid6               (hip_pipe_rxvalid6), //                   .rxvalid6
		.rxvalid7               (hip_pipe_rxvalid7), //                   .rxvalid7
		.app_int_sts            (apps_int_msi_app_int_sts),  //            int_msi.app_int_sts
		.app_msi_num            (apps_int_msi_app_msi_num),  //                   .app_msi_num
		.app_msi_req            (apps_int_msi_app_msi_req),  //                   .app_msi_req
		.app_msi_tc             (apps_int_msi_app_msi_tc),   //                   .app_msi_tc
		.app_int_ack            (pcie_gen2x8_inst_int_msi_app_int_ack),  //                   .app_int_ack
		.app_msi_ack            (pcie_gen2x8_inst_int_msi_app_msi_ack),  //                   .app_msi_ack
		.test_in                (iHIP_CTRL_TEST_IN),  //           hip_ctrl.test_in
		.simu_mode_pipe         (iHIP_CTRL_SIMU_MODE_PIPE),   //                   .simu_mode_pipe
		.derr_cor_ext_rcv       (pcie_gen2x8_inst_hip_status_derr_cor_ext_rcv),  //         hip_status.derr_cor_ext_rcv
		.derr_cor_ext_rpl       (pcie_gen2x8_inst_hip_status_derr_cor_ext_rpl),  //                   .derr_cor_ext_rpl
		.derr_rpl               (pcie_gen2x8_inst_hip_status_derr_rpl),  //                   .derr_rpl
		.dlup                   (pcie_gen2x8_inst_hip_status_dlup),      //                   .dlup
		.dlup_exit              (pcie_gen2x8_inst_hip_status_dlup_exit), //                   .dlup_exit
		.ev128ns                (pcie_gen2x8_inst_hip_status_ev128ns),   //                   .ev128ns
		.ev1us                  (pcie_gen2x8_inst_hip_status_ev1us),     //                   .ev1us
		.hotrst_exit            (pcie_gen2x8_inst_hip_status_hotrst_exit),       //                   .hotrst_exit
		.int_status             (pcie_gen2x8_inst_hip_status_int_status),//                   .int_status
		.l2_exit                (pcie_gen2x8_inst_hip_status_l2_exit),   //                   .l2_exit
		.lane_act               (pcie_gen2x8_inst_hip_status_lane_act),  //                   .lane_act
		.ltssmstate             (pcie_gen2x8_inst_hip_status_ltssmstate),//                   .ltssmstate
		.rx_par_err             (pcie_gen2x8_inst_hip_status_rx_par_err),//                   .rx_par_err
		.tx_par_err             (pcie_gen2x8_inst_hip_status_tx_par_err),//                   .tx_par_err
		.cfg_par_err            (pcie_gen2x8_inst_hip_status_cfg_par_err),       //                   .cfg_par_err
		.ko_cpl_spc_header      (pcie_gen2x8_inst_hip_status_ko_cpl_spc_header), //                   .ko_cpl_spc_header
		.ko_cpl_spc_data        (pcie_gen2x8_inst_hip_status_ko_cpl_spc_data),   //                   .ko_cpl_spc_data
		.currentspeed           (pcie_gen2x8_inst_hip_currentspeed_currentspeed),//   hip_currentspeed.currentspeed
		.rx_st_parity           (),                  //        (terminated)
		.tx_st_parity           (32'b00000000000000000000000000000000),  //        (terminated)
		.tx_cons_cred_sel       (1'b0),              //        (terminated)
		.sim_pipe_pclk_out      (),                  //        (terminated)
		.rxdataskip0            (1'b0),              //        (terminated)
		.rxdataskip1            (1'b0),              //        (terminated)
		.rxdataskip2            (1'b0),              //        (terminated)
		.rxdataskip3            (1'b0),              //        (terminated)
		.rxdataskip4            (1'b0),              //        (terminated)
		.rxdataskip5            (1'b0),              //        (terminated)
		.rxdataskip6            (1'b0),              //        (terminated)
		.rxdataskip7            (1'b0),              //        (terminated)
		.rxblkst0               (1'b0),              //        (terminated)
		.rxblkst1               (1'b0),              //        (terminated)
		.rxblkst2               (1'b0),              //        (terminated)
		.rxblkst3               (1'b0),              //        (terminated)
		.rxblkst4               (1'b0),              //        (terminated)
		.rxblkst5               (1'b0),              //        (terminated)
		.rxblkst6               (1'b0),              //        (terminated)
		.rxblkst7               (1'b0),              //        (terminated)
		.rxsynchd0              (2'b00),             //        (terminated)
		.rxsynchd1              (2'b00),             //        (terminated)
		.rxsynchd2              (2'b00),             //        (terminated)
		.rxsynchd3              (2'b00),             //        (terminated)
		.rxsynchd4              (2'b00),             //        (terminated)
		.rxsynchd5              (2'b00),             //        (terminated)
		.rxsynchd6              (2'b00),             //        (terminated)
		.rxsynchd7              (2'b00),             //        (terminated)
		.rxfreqlocked0          (1'b0),              //        (terminated)
		.rxfreqlocked1          (1'b0),              //        (terminated)
		.rxfreqlocked2          (1'b0),              //        (terminated)
		.rxfreqlocked3          (1'b0),              //        (terminated)
		.rxfreqlocked4          (1'b0),              //        (terminated)
		.rxfreqlocked5          (1'b0),              //        (terminated)
		.rxfreqlocked6          (1'b0),              //        (terminated)
		.rxfreqlocked7          (1'b0),              //        (terminated)
		.currentcoeff0          (),                  //        (terminated)
		.currentcoeff1          (),                  //        (terminated)
		.currentcoeff2          (),                  //        (terminated)
		.currentcoeff3          (),                  //        (terminated)
		.currentcoeff4          (),                  //        (terminated)
		.currentcoeff5          (),                  //        (terminated)
		.currentcoeff6          (),                  //        (terminated)
		.currentcoeff7          (),                  //        (terminated)
		.currentrxpreset0       (),                  //        (terminated)
		.currentrxpreset1       (),                  //        (terminated)
		.currentrxpreset2       (),                  //        (terminated)
		.currentrxpreset3       (),                  //        (terminated)
		.currentrxpreset4       (),                  //        (terminated)
		.currentrxpreset5       (),                  //        (terminated)
		.currentrxpreset6       (),                  //        (terminated)
		.currentrxpreset7       (),                  //        (terminated)
		.txsynchd0              (),                  //        (terminated)
		.txsynchd1              (),                  //        (terminated)
		.txsynchd2              (),                  //        (terminated)
		.txsynchd3              (),                  //        (terminated)
		.txsynchd4              (),                  //        (terminated)
		.txsynchd5              (),                  //        (terminated)
		.txsynchd6              (),                  //        (terminated)
		.txsynchd7              (),                  //        (terminated)
		.txblkst0               (),                  //        (terminated)
		.txblkst1               (),                  //        (terminated)
		.txblkst2               (),                  //        (terminated)
		.txblkst3               (),                  //        (terminated)
		.txblkst4               (),                  //        (terminated)
		.txblkst5               (),                  //        (terminated)
		.txblkst6               (),                  //        (terminated)
		.txblkst7               (),                  //        (terminated)
		.aer_msi_num            (5'b00000),          //        (terminated)
		.pex_msi_num            (5'b00000),          //        (terminated)
		.serr_out               (),                  //        (terminated)
		.hip_reconfig_clk       (1'b0),              //        (terminated)
		.hip_reconfig_rst_n     (1'b0),              //        (terminated)
		.hip_reconfig_address   (10'b0000000000),    //        (terminated)
		.hip_reconfig_read      (1'b0),              //        (terminated)
		.hip_reconfig_write     (1'b0),              //        (terminated)
		.hip_reconfig_writedata (16'b0000000000000000),      //        (terminated)
		.hip_reconfig_byte_en   (2'b00),             //        (terminated)
		.ser_shift_load         (1'b0),              //        (terminated)
		.interface_sel          (1'b0),              //        (terminated)
		.cfgbp_link2csr         (13'b0000000000000), //        (terminated)
		.cfgbp_comclk_reg       (1'b0),              //        (terminated)
		.cfgbp_extsy_reg        (1'b0),              //        (terminated)
		.cfgbp_max_pload        (3'b000),            //        (terminated)
		.cfgbp_tx_ecrcgen       (1'b0),              //        (terminated)
		.cfgbp_rx_ecrchk        (1'b0),              //        (terminated)
		.cfgbp_secbus           (8'b00000000),       //        (terminated)
		.cfgbp_linkcsr_bit0     (1'b0),              //        (terminated)
		.cfgbp_tx_req_pm        (1'b0),              //        (terminated)
		.cfgbp_tx_typ_pm        (3'b000),            //        (terminated)
		.cfgbp_req_phypm        (4'b0000),           //        (terminated)
		.cfgbp_req_phycfg       (4'b0000),           //        (terminated)
		.cfgbp_vc0_tcmap_pld    (7'b0000000),        //        (terminated)
		.cfgbp_inh_dllp         (1'b0),              //        (terminated)
		.cfgbp_inh_tx_tlp       (1'b0),              //        (terminated)
		.cfgbp_req_wake         (1'b0),              //        (terminated)
		.cfgbp_link3_ctl        (2'b00),             //        (terminated)
		.cseb_rddata            (32'b00000000000000000000000000000000),  //        (terminated)
		.cseb_rdresponse        (5'b00000),          //        (terminated)
		.cseb_waitrequest       (1'b0),              //        (terminated)
		.cseb_wrresponse        (5'b00000),          //        (terminated)
		.cseb_wrresp_valid      (1'b0),              //        (terminated)
		.cseb_rddata_parity     (4'b0000),           //        (terminated)
		.reservedin             (32'b00000000000000000000000000000000),  //        (terminated)
		.tlbfm_in               (),                  //        (terminated)
		.tlbfm_out              (1001'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000), //        (terminated)
		.rxfc_cplbuf_ovf        ()                   //        (terminated)
	);

`ifdef NOHIP
assign apps_tx_st_data  = 256'h0;   
assign apps_tx_st_empty = 2'h1;  
assign apps_tx_st_endofpacket   = 1'b0;    
assign apps_tx_st_error   = 1'b0;    
assign apps_tx_st_startofpacket   = 1'b0;    
assign apps_tx_st_valid = 1'b0;     
`endif   

bali_pcie_app #(
    .PORTS      ( PORTS             ),
    .BALI       ( BALI              )
)
bali_pcie_app_inst
(
    .tx_cred_datafccp       (pcie_gen2x8_inst_tx_cred_tx_cred_datafccp),     //            tx_cred.tx_cred_datafccp
    .tx_cred_datafcnp       (pcie_gen2x8_inst_tx_cred_tx_cred_datafcnp),     //                   .tx_cred_datafcnp
    .tx_cred_datafcp        (pcie_gen2x8_inst_tx_cred_tx_cred_datafcp),      //                   .tx_cred_datafcp
    .tx_cred_fchipcons      (pcie_gen2x8_inst_tx_cred_tx_cred_fchipcons),    //                   .tx_cred_fchipcons
    .tx_cred_fcinfinite     (pcie_gen2x8_inst_tx_cred_tx_cred_fcinfinite),   //                   .tx_cred_fcinfinite
    .tx_cred_hdrfccp        (pcie_gen2x8_inst_tx_cred_tx_cred_hdrfccp),      //                   .tx_cred_hdrfccp
    .tx_cred_hdrfcnp        (pcie_gen2x8_inst_tx_cred_tx_cred_hdrfcnp),      //                   .tx_cred_hdrfcnp
    .tx_cred_hdrfcp         (pcie_gen2x8_inst_tx_cred_tx_cred_hdrfcp),       //                   .tx_cred_hdrfcp

  //////////////////////////////////////////////////////////////////////
  // TO/FROM TOP-LEVEL MM REG DECODE I/F
  //////////////////////////////////////////////////////////////////////
 .oPCIE2MM_WR_DATA        (oPCIE2MM_WR_DATA),
 .oPCIE2MM_ADDRESS        (oPCIE2MM_ADDRESS),
 .oPCIE2MM_WR_EN          (oPCIE2MM_WR_EN),
 .oPCIE2MM_RD_EN          (oPCIE2MM_RD_EN),
 .iMM2PCIE_ACK            (iMM2PCIE_ACK),
 .iMM2PCIE_RD_DATA        (iMM2PCIE_RD_DATA),
  //////////////////////////////////////////////////////////////////////
  // TO/FROM MM REG DECODE I/F
  //////////////////////////////////////////////////////////////////////
  .iMM_WR_DATA            (iMM_WR_DATA),
  .iMM_ADDR               (iMM_ADDR),
  .iMM_WR_EN              (iMM_WR_EN),
  .iMM_RD_EN              (iMM_RD_EN),
  .oMM_RD_DATA            (oMM_RD_DATA),
  .oMM_RD_DATA_V          (oMM_RD_DATA_V),

  //////////////////////////////////////////////////////////////////////
  // DMA WRITE to DPL BUFFER I/F
  //////////////////////////////////////////////////////////////////////
  .iDPLBUF_REQ           (iDPLBUF_REQ),
  .oDPLBUF_GNT           (oDPLBUF_GNT),
  .iDPLBUF_DATA          (iDPLBUF_DATA),
  .iDPLBUF_DATA_V        (iDPLBUF_DATA_V),

  .oAPP_RST_n_STATUS     (oAPP_RST_n_STATUS),

`ifdef NOHIP
 .oTX_ST_DATA                           (),     // 
 .oTX_ST_EMPTY                          (),      // 
 .oTX_ST_EOP                            (),             // 
 .oTX_ST_ERR                            (),             // 
 .oTX_ST_SOP                            (),             // 
 .oTX_ST_VALID                          (),           // 
 //.oTX_ST_PARITY                         (apps_tx_st_parity[31:0]),    // <<< NOT USED
 .iTX_ST_READY                          (),           // 
`else
 .oTX_ST_DATA                           (apps_tx_st_data[255:0]),     // 
 .oTX_ST_EMPTY                          (apps_tx_st_empty[1:0]),      // 
 .oTX_ST_EOP                            (apps_tx_st_endofpacket),             // 
 .oTX_ST_ERR                            (apps_tx_st_error),             // 
 .oTX_ST_SOP                            (apps_tx_st_startofpacket),             // 
 .oTX_ST_VALID                          (apps_tx_st_valid),           // 
 //.oTX_ST_PARITY                         (apps_tx_st_parity[31:0]),    // <<< NOT USED
 .iTX_ST_READY                          (apps_tx_st_ready),           // 
`endif
 
 .iCLK_PCIE_CORECLKOUT_HIP              (oCLK_PCIE_CORECLKOUT_HIP),
 /*AUTOINST*/
 // Outputs
.oA2HIP_PLD_CORE_READY                 (apps_hip_rst_pld_core_ready),  // 
 //.oA2HIP_RECONFIG_TO_XCVR               (a2hip_reconfig_to_xcvr[700-1:0]), // <<<REMOVE, extern reconfig
 //.oA2HIP_BUSY_XCVR_RECONFIG             (a2hip_busy_xcvr_reconfig), // <<<REMOVE, extern reconfig
 .oA2HIP_LMI_ADDR                       (apps_lmi_lmi_addr),  // 
 .oA2HIP_LMI_DIN                        (apps_lmi_lmi_din[31:0]),   // 
 .oA2HIP_LMI_RDEN                       (apps_lmi_lmi_rden),        // 
 .oA2HIP_LMI_WREN                       (apps_lmi_lmi_wren),        // 
 .oA2HIP_PM_AUXPWR                      (apps_power_mngt_pm_auxpwr),       // 
 .oA2HIP_PM_DATA                        (apps_power_mngt_pm_data[9:0]),    // 
 .oA2HIP_PME_TO_CR                      (apps_power_mngt_pme_to_cr),       // 
 .oA2HIP_PM_EVENT                       (apps_power_mngt_pm_event),        // 
 //.oA2HIP_PM_EVENT_FUNC                  (a2hip_pm_event_func[2:0]), // <<< NOT USED
 .oRX_ST_READY                          (pcie_gen2x8_inst_rx_st_ready),           // 
 .oRX_ST_MASK                           (apps_rx_bar_be_rx_st_mask),            // 
 //.oCFGLINK2CSRPLD                       (cfglink2csrpld[12:0]),  // <<< NOT USED
 .oA2HIP_CPL_ERR                        (apps_config_tl_cpl_err),    // 
 .oA2HIP_CPL_PENDING                    (apps_config_tl_cpl_pending),     // 
 //.oA2HIP_CPL_ERR_FUNC                   (a2hip_cpl_err_func[2:0]), // <<< NOT USED
 // Inputs
 .iHIP2A_RESET_STATUS                   (pcie_gen2x8_inst_hip_rst_reset_status),    // 
 .iHIP2A_SERDES_PLL_LOCKED              (pcie_gen2x8_inst_hip_rst_serdes_pll_locked), // 
 .iHIP2A_PLD_CLK_INUSE                  (pcie_gen2x8_inst_hip_rst_pld_clk_inuse),   // 
 .iCLK_PCIE_GLOBAL                      (iCLK_PCIE_GLOBAL),      // 
 .testin_zero                           (pcie_gen2x8_inst_hip_rst_testin_zero),          //     <<<ADD NEW
                .app_int_sts            (apps_int_msi_app_int_sts),  //            int_msi.app_int_sts  <<<ADD NEW, drive 0
                .app_msi_num            (apps_int_msi_app_msi_num),  //                   .app_msi_num  <<<ADD NEW, drive 0
                .app_msi_req            (apps_int_msi_app_msi_req),  //                   .app_msi_req  <<<ADD NEW, drive 0
                .app_msi_tc             (apps_int_msi_app_msi_tc),   //                   .app_msi_tc  <<<ADD NEW, drive 0
                .app_int_ack            (pcie_gen2x8_inst_int_msi_app_int_ack),  //                   .app_int_ack  <<<ADD NEW, expect 0
                .app_msi_ack            (pcie_gen2x8_inst_int_msi_app_msi_ack),  //                   .app_msi_ack  <<<ADD NEW, expect 0

                .derr_cor_ext_rcv_drv  (apps_hip_status_drv_derr_cor_ext_rcv),          // hip_status_drv.derr_cor_ext_rcv  <<<ADD NEW, flop then drive 
                .derr_cor_ext_rpl_drv  (apps_hip_status_drv_derr_cor_ext_rpl),          //               .derr_cor_ext_rpl  <<<ADD NEW, flop then drive 
                .derr_rpl_drv          (apps_hip_status_drv_derr_rpl),                  //               .derr_rpl  <<<ADD NEW, flop then drive 
                .dlup_exit_drv         (apps_hip_status_drv_dlup_exit),                 //               .dlup_exit  <<<ADD NEW, flop then drive 
                .ev128ns_drv           (apps_hip_status_drv_ev128ns),                   //               .ev128ns  <<<ADD NEW, flop then drive 
                .ev1us_drv             (apps_hip_status_drv_ev1us),                     //               .ev1us  <<<ADD NEW, flop then drive 
                .hotrst_exit_drv       (apps_hip_status_drv_hotrst_exit),               //               .hotrst_exit  <<<ADD NEW, flop then drive 
                .int_status_drv        (apps_hip_status_drv_int_status),                //               .int_status  <<<ADD NEW, flop then drive 
                .l2_exit_drv           (apps_hip_status_drv_l2_exit),                   //               .l2_exit  <<<ADD NEW, flop then drive 
                .lane_act_drv          (apps_hip_status_drv_lane_act),                  //               .lane_act  <<<ADD NEW, flop then drive 
                .ltssmstate_drv        (apps_hip_status_drv_ltssmstate),                //               .ltssmstate  <<<ADD NEW, flop then drive 
                .dlup_drv              (apps_hip_status_drv_dlup),                      //               .dlup  <<<ADD NEW, flop then drive 
                .rx_par_err_drv        (apps_hip_status_drv_rx_par_err),                //               .rx_par_err  <<<ADD NEW, flop then drive 
                .tx_par_err_drv        (apps_hip_status_drv_tx_par_err),                //               .tx_par_err  <<<ADD NEW, flop then drive 
                .cfg_par_err_drv       (apps_hip_status_drv_cfg_par_err),               //               .cfg_par_err  <<<ADD NEW, flop then drive 
                .ko_cpl_spc_header_drv (apps_hip_status_drv_ko_cpl_spc_header),         //               .ko_cpl_spc_header  <<<ADD NEW, flop then drive 
                .ko_cpl_spc_data_drv   (apps_hip_status_drv_ko_cpl_spc_data),           //               .ko_cpl_spc_data  <<<ADD NEW, flop then drive 
                .hpg_ctrler            (apps_config_tl_hpg_ctrler),                     //      config_tl.hpg_ctrler  <<<ADD NEW, drive 0


 .iRST_100M_N                           (iRST_100M_N),           // Templated
 .iRST_PCIE_N                           (iRST_PCIE_N),           // Templated
 .iRST_CHIP_PCIE_N                      (iRST_CHIP_PCIE_N),           // Templated
 .iCLK_100M                             (iCLK_100M),             // 
 .iRECONFIG_XCVR_CLK                    (iRECONFIG_XCVR_CLK),     // 
 //.iHIP2APP_RECONFIG_FROM_XCVR           (hip2app_reconfig_from_xcvr[459:0]), // <<<REMOVE, extern reconfig
 .iHIP2A_TL_CFG_ADD                     (pcie_gen2x8_inst_config_tl_tl_cfg_add), // 
 .iHIP2A_TL_CFG_CTL                     (pcie_gen2x8_inst_config_tl_tl_cfg_ctl), // 
 .iHIP2A_TL_CFG_STS                     (pcie_gen2x8_inst_config_tl_tl_cfg_sts), // 
 .iHIP2A_LMI_ACK                        (pcie_gen2x8_inst_lmi_lmi_ack),         // 
 .iHIP2A_LMI_DOUT                       (pcie_gen2x8_inst_lmi_lmi_dout),  // 
 .iHIP2A_PME_TO_SR                      (pcie_gen2x8_inst_power_mngt_pme_to_sr),       // 
 .iRX_ST_DATA                           (pcie_gen2x8_inst_rx_st_data),     // 
 .iRX_ST_SOP                            (pcie_gen2x8_inst_rx_st_startofpacket),             // 
 .iRX_ST_VALID                          (pcie_gen2x8_inst_rx_st_valid),           // 
 .iRX_ST_EMPTY                          (pcie_gen2x8_inst_rx_st_empty),      // 
 .iRX_ST_EOP                            (pcie_gen2x8_inst_rx_st_endofpacket),             // 
 .iRX_ST_ERR                            (pcie_gen2x8_inst_rx_st_error),             // 
 .iRX_ST_BE                             (pcie_gen2x8_inst_rx_bar_be_rx_st_be),        // 
 .iRX_ST_BAR                            (pcie_gen2x8_inst_rx_bar_be_rx_st_bar),        // 
 .iHIP2A_CURRENTSPEED                   (pcie_gen2x8_inst_hip_currentspeed_currentspeed), // 
 .iHIP2A_DERR_COR_EXT_RCV               (pcie_gen2x8_inst_hip_status_derr_cor_ext_rcv), // 
 .iHIP2A_DERR_COR_EXT_RPL               (pcie_gen2x8_inst_hip_status_derr_cor_ext_rpl), // 
 .iHIP2A_DERR_RPL                       (pcie_gen2x8_inst_hip_status_derr_rpl),        // 
 .iHIP2A_RX_PAR_ERR                     (pcie_gen2x8_inst_hip_status_rx_par_err),      // 
 .iHIP2A_TX_PAR_ERR                     (pcie_gen2x8_inst_hip_status_tx_par_err), // 
 .iHIP2A_CFG_PAR_ERR                    (pcie_gen2x8_inst_hip_status_cfg_par_err),     // 
 .iHIP2A_DLUP                           (pcie_gen2x8_inst_hip_status_dlup),            // 
 .iHIP2A_DLUP_EXIT_n                    (pcie_gen2x8_inst_hip_status_dlup_exit),     // 
 .iHIP2A_EV128NS                        (pcie_gen2x8_inst_hip_status_ev128ns),         // 
 .iHIP2A_EV1US                          (pcie_gen2x8_inst_hip_status_ev1us),           // 
 .iHIP2A_HOTRST_EXIT_n                  (pcie_gen2x8_inst_hip_status_hotrst_exit),   // 
 .iHIP2A_INT_STATUS                     (pcie_gen2x8_inst_hip_status_int_status), // 
 .iHIP2A_L2_EXIT_n                      (pcie_gen2x8_inst_hip_status_l2_exit),       // 
 .iHIP2A_LANE_ACT                       (pcie_gen2x8_inst_hip_status_lane_act),   // 
 .iHIP2A_LTSSMSTATE                     (pcie_gen2x8_inst_hip_status_ltssmstate), // 
 .iHIP2A_KO_CPL_SPC_HEADER              (pcie_gen2x8_inst_hip_status_ko_cpl_spc_header), //
 .iHIP2A_KO_CPL_SPC_DATA                (pcie_gen2x8_inst_hip_status_ko_cpl_spc_data)
);

	altpcie_reconfig_driver #(
		.INTENDED_DEVICE_FAMILY        ("Stratix V"),
		.gen123_lane_rate_mode_hwtcl   ("Gen2 (5.0 Gbps)"),
		.number_of_reconfig_interfaces (11)
	) pcie_reconfig_driver_0 (
		.reconfig_xcvr_clk         (iRECONFIG_XCVR_CLK),                                          // reconfig_xcvr_clk.clk
		.reconfig_xcvr_rst         (rst_controller_reset_out_reset),                   // reconfig_xcvr_rst.reset
		.reconfig_mgmt_address     (pcie_reconfig_driver_0_reconfig_mgmt_address),     //     reconfig_mgmt.address
		.reconfig_mgmt_read        (pcie_reconfig_driver_0_reconfig_mgmt_read),        //                  .read
		.reconfig_mgmt_readdata    (pcie_reconfig_driver_0_reconfig_mgmt_readdata),    //                  .readdata
		.reconfig_mgmt_waitrequest (pcie_reconfig_driver_0_reconfig_mgmt_waitrequest), //                  .waitrequest
		.reconfig_mgmt_write       (pcie_reconfig_driver_0_reconfig_mgmt_write),       //                  .write
		.reconfig_mgmt_writedata   (pcie_reconfig_driver_0_reconfig_mgmt_writedata),   //                  .writedata
		.currentspeed              (pcie_gen2x8_inst_hip_currentspeed_currentspeed),   //  hip_currentspeed.currentspeed
		.reconfig_busy             (alt_xcvr_reconfig_0_reconfig_busy_reconfig_busy),  //     reconfig_busy.reconfig_busy
		.pld_clk                   (iCLK_PCIE_GLOBAL),                             //           pld_clk.clk
		.derr_cor_ext_rcv_drv      (apps_hip_status_drv_derr_cor_ext_rcv),             //    hip_status_drv.derr_cor_ext_rcv
		.derr_cor_ext_rpl_drv      (apps_hip_status_drv_derr_cor_ext_rpl),             //                  .derr_cor_ext_rpl
		.derr_rpl_drv              (apps_hip_status_drv_derr_rpl),                     //                  .derr_rpl
		.dlup_exit_drv             (apps_hip_status_drv_dlup_exit),                    //                  .dlup_exit
		.ev128ns_drv               (apps_hip_status_drv_ev128ns),                      //                  .ev128ns
		.ev1us_drv                 (apps_hip_status_drv_ev1us),                        //                  .ev1us
		.hotrst_exit_drv           (apps_hip_status_drv_hotrst_exit),                  //                  .hotrst_exit
		.int_status_drv            (apps_hip_status_drv_int_status),                   //                  .int_status
		.l2_exit_drv               (apps_hip_status_drv_l2_exit),                      //                  .l2_exit
		.lane_act_drv              (apps_hip_status_drv_lane_act),                     //                  .lane_act
		.ltssmstate_drv            (apps_hip_status_drv_ltssmstate),                   //                  .ltssmstate
		.dlup_drv                  (apps_hip_status_drv_dlup),                         //                  .dlup
		.rx_par_err_drv            (apps_hip_status_drv_rx_par_err),                   //                  .rx_par_err
		.tx_par_err_drv            (apps_hip_status_drv_tx_par_err),                   //                  .tx_par_err
		.cfg_par_err_drv           (apps_hip_status_drv_cfg_par_err),                  //                  .cfg_par_err
		.ko_cpl_spc_header_drv     (apps_hip_status_drv_ko_cpl_spc_header),            //                  .ko_cpl_spc_header
		.ko_cpl_spc_data_drv       (apps_hip_status_drv_ko_cpl_spc_data),              //                  .ko_cpl_spc_data
		.cal_busy_in               ()                                                  //       (terminated)
	);

generate 
  if (BALI == 1) begin : gen_extr_reconf
  alt_xcvr_reconfig #(
    .device_family                 ("Stratix V"),
    .number_of_reconfig_interfaces (12),
    .enable_offset                 (1),
    .enable_lc                     (1),
    .enable_dcd                    (0),
    .enable_dcd_power_up           (1),
    .enable_analog                 (0),
    .enable_eyemon                 (0),
    .enable_ber                    (0),
    .enable_dfe                    (0),
    .enable_adce                   (0),
    .enable_mif                    (0),
    .enable_pll                    (0)
  ) alt_xcvr_reconfig_0 (
    .reconfig_busy             (alt_xcvr_reconfig_0_reconfig_busy_reconfig_busy),        //      reconfig_busy.reconfig_busy
    .mgmt_clk_clk              (iRECONFIG_XCVR_CLK),                                                //       mgmt_clk_clk.clk
    .mgmt_rst_reset            (rst_controller_reset_out_reset),                         //     mgmt_rst_reset.reset
    .reconfig_mgmt_address     (pcie_reconfig_driver_0_reconfig_mgmt_address),           //      reconfig_mgmt.address
    .reconfig_mgmt_read        (pcie_reconfig_driver_0_reconfig_mgmt_read),              //                   .read
    .reconfig_mgmt_readdata    (pcie_reconfig_driver_0_reconfig_mgmt_readdata),          //                   .readdata
    .reconfig_mgmt_waitrequest (pcie_reconfig_driver_0_reconfig_mgmt_waitrequest),       //                   .waitrequest
    .reconfig_mgmt_write       (pcie_reconfig_driver_0_reconfig_mgmt_write),             //                   .write
    .reconfig_mgmt_writedata   (pcie_reconfig_driver_0_reconfig_mgmt_writedata),         //                   .writedata
    .reconfig_to_xcvr          ({fc_reconfig_to_xcvr, alt_xcvr_reconfig_0_reconfig_to_xcvr_reconfig_to_xcvr}),  //   reconfig_to_xcvr.reconfig_to_xcvr
    .reconfig_from_xcvr        ({fc_reconfig_from_xcvr, pcie_gen2x8_inst_reconfig_from_xcvr_reconfig_from_xcvr}), // reconfig_from_xcvr.reconfig_from_xcvr
    .tx_cal_busy               (),                                                       //        (terminated)
    .rx_cal_busy               (),                                                       //        (terminated)
    .cal_busy_in               (1'b0),                                                   //        (terminated)
    .reconfig_mif_address      (),                                                       //        (terminated)
    .reconfig_mif_read         (),                                                       //        (terminated)
    .reconfig_mif_readdata     (16'b0000000000000000),                                   //        (terminated)
    .reconfig_mif_waitrequest  (1'b0)                                                    //        (terminated)
  );

	end : gen_extr_reconf

  else begin : gen_normal 
	alt_xcvr_reconfig #(
		.device_family                 ("Stratix V"),
		.number_of_reconfig_interfaces (11),
		.enable_offset                 (1),
		.enable_lc                     (1),
		.enable_dcd                    (0),
		.enable_dcd_power_up           (1),
		.enable_analog                 (0),
		.enable_eyemon                 (0),
		.enable_ber                    (0),
		.enable_dfe                    (0),
		.enable_adce                   (0),
		.enable_mif                    (0),
		.enable_pll                    (0)
	) alt_xcvr_reconfig_0 (
		.reconfig_busy             (alt_xcvr_reconfig_0_reconfig_busy_reconfig_busy),        //      reconfig_busy.reconfig_busy
		.mgmt_clk_clk              (iRECONFIG_XCVR_CLK),                                                //       mgmt_clk_clk.clk
		.mgmt_rst_reset            (rst_controller_reset_out_reset),                         //     mgmt_rst_reset.reset
		.reconfig_mgmt_address     (pcie_reconfig_driver_0_reconfig_mgmt_address),           //      reconfig_mgmt.address
		.reconfig_mgmt_read        (pcie_reconfig_driver_0_reconfig_mgmt_read),              //                   .read
		.reconfig_mgmt_readdata    (pcie_reconfig_driver_0_reconfig_mgmt_readdata),          //                   .readdata
		.reconfig_mgmt_waitrequest (pcie_reconfig_driver_0_reconfig_mgmt_waitrequest),       //                   .waitrequest
		.reconfig_mgmt_write       (pcie_reconfig_driver_0_reconfig_mgmt_write),             //                   .write
		.reconfig_mgmt_writedata   (pcie_reconfig_driver_0_reconfig_mgmt_writedata),         //                   .writedata
		.reconfig_to_xcvr          (alt_xcvr_reconfig_0_reconfig_to_xcvr_reconfig_to_xcvr),  //   reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr        (pcie_gen2x8_inst_reconfig_from_xcvr_reconfig_from_xcvr), // reconfig_from_xcvr.reconfig_from_xcvr
		.tx_cal_busy               (),                                                       //        (terminated)
		.rx_cal_busy               (),                                                       //        (terminated)
		.cal_busy_in               (1'b0),                                                   //        (terminated)
		.reconfig_mif_address      (),                                                       //        (terminated)
		.reconfig_mif_read         (),                                                       //        (terminated)
		.reconfig_mif_readdata     (16'b0000000000000000),                                   //        (terminated)
		.reconfig_mif_waitrequest  (1'b0)                                                    //        (terminated)
	);
  end : gen_normal
endgenerate

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		//lz change sync method .OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.OUTPUT_RESET_SYNC_EDGES ("none"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		//lz try different reset .reset_in0  (~iRST_NPOR_n),                 // reset_in0.reset
		.reset_in0  (~iPIN_PERST_n),                 // reset_in0.reset
		.clk        (iRECONFIG_XCVR_CLK),                        //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

 assign oLANE_ACT = pcie_gen2x8_inst_hip_status_lane_act;
 assign oLTSSM    = pcie_gen2x8_inst_hip_status_ltssmstate;
 assign oCURRENT_SPEED = pcie_gen2x8_inst_hip_currentspeed_currentspeed;

reg heart_beat;

always @ (posedge iRECONFIG_XCVR_CLK or negedge iPIN_PERST_n)
  if (!iPIN_PERST_n)
    heart_beat <= 1'b1;
  else
    heart_beat <= !heart_beat;

assign oPCIE_MISC_STATUS =
                            {7'h0,
                             heart_beat,
                             iRST_NPOR_n,
                             pcie_gen2x8_inst_hip_status_lane_act,
                             pcie_gen2x8_inst_hip_currentspeed_currentspeed,
                             rst_controller_reset_out_reset,
                             oLTSSM,
                             oAPP_RST_n_STATUS,
                             pcie_gen2x8_inst_hip_status_dlup_exit,           // 1 - pulses 1-0-1 on exit from data link up
                             pcie_gen2x8_inst_hip_status_hotrst_exit,         // 1 - pulses 1-0-1

                             pcie_gen2x8_inst_hip_status_l2_exit,              //1 -> pulses 1-0-1 to tell app to reset for 32 cycles
                             pcie_gen2x8_inst_hip_status_dlup,                  // 1 - good
                             alt_xcvr_reconfig_0_reconfig_busy_reconfig_busy,    // 0 - good
                             pcie_gen2x8_inst_hip_rst_reset_status,          // 0 - good - reset sequence shows going 1 to 0, then holding 0 if 32-cycles between de-assert of pld_clk_inuse to deassert of crst/srst

                             pcie_gen2x8_inst_hip_rst_serdes_pll_locked,     // 1 - good
                             apps_hip_rst_pld_core_ready,        // 1 - good
                             pcie_gen2x8_inst_hip_rst_pld_clk_inuse,         // 1 - good
                             iPIN_PERST_n                 // 1 - MB not resetting PCIE
                             };

//signaltap signal_tap_inst(
        //.acq_clk(iRECONFIG_XCVR_CLK),
        //.acq_data_in(oPCIE_MISC_STATUS),
        //.acq_trigger_in({3'h0, oLTSSM})
//);

endmodule
